
module FD_0 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_96 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_95 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_94 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_93 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_92 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_91 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_90 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_89 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_88 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_87 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_86 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_85 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_84 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_83 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_82 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_81 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_80 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_79 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_78 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_77 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_76 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_75 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_74 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_73 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_72 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_71 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_70 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_69 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_68 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_67 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_66 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_GENERIC_NBIT32_0 ( D, CLK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET;
  wire   n1, n2, n3;

  FD_0 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n3), .Q(Q[0]) );
  FD_96 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n1), .Q(Q[1]) );
  FD_95 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n1), .Q(Q[2]) );
  FD_94 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n1), .Q(Q[3]) );
  FD_93 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n1), .Q(Q[4]) );
  FD_92 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n1), .Q(Q[5]) );
  FD_91 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n1), .Q(Q[6]) );
  FD_90 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n1), .Q(Q[7]) );
  FD_89 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n1), .Q(Q[8]) );
  FD_88 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n1), .Q(Q[9]) );
  FD_87 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n1), .Q(Q[10]) );
  FD_86 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n1), .Q(Q[11]) );
  FD_85 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n1), .Q(Q[12]) );
  FD_84 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n2), .Q(Q[13]) );
  FD_83 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n2), .Q(Q[14]) );
  FD_82 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n2), .Q(Q[15]) );
  FD_81 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n2), .Q(Q[16]) );
  FD_80 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n2), .Q(Q[17]) );
  FD_79 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n2), .Q(Q[18]) );
  FD_78 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n2), .Q(Q[19]) );
  FD_77 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n2), .Q(Q[20]) );
  FD_76 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n2), .Q(Q[21]) );
  FD_75 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n2), .Q(Q[22]) );
  FD_74 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n2), .Q(Q[23]) );
  FD_73 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n2), .Q(Q[24]) );
  FD_72 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n3), .Q(Q[25]) );
  FD_71 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n3), .Q(Q[26]) );
  FD_70 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n3), .Q(Q[27]) );
  FD_69 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n3), .Q(Q[28]) );
  FD_68 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n3), .Q(Q[29]) );
  FD_67 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n3), .Q(Q[30]) );
  FD_66 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n1) );
  BUF_X1 U2 ( .A(RESET), .Z(n2) );
  BUF_X1 U3 ( .A(RESET), .Z(n3) );
endmodule


module FD_65 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_64 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_63 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_62 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_61 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_60 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_59 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_58 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_57 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_56 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_55 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_54 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_53 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_52 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_51 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_50 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_49 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_48 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_47 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_46 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_45 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_44 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_43 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_42 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_41 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_40 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_39 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_38 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_37 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_36 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_35 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_34 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_GENERIC_NBIT32_1 ( D, CLK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET;
  wire   n1, n2, n3;

  FD_65 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n1), .Q(Q[0]) );
  FD_64 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n1), .Q(Q[1]) );
  FD_63 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n1), .Q(Q[2]) );
  FD_62 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n1), .Q(Q[3]) );
  FD_61 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n1), .Q(Q[4]) );
  FD_60 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n1), .Q(Q[5]) );
  FD_59 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n1), .Q(Q[6]) );
  FD_58 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n1), .Q(Q[7]) );
  FD_57 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n1), .Q(Q[8]) );
  FD_56 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n1), .Q(Q[9]) );
  FD_55 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n1), .Q(Q[10]) );
  FD_54 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n1), .Q(Q[11]) );
  FD_53 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n2), .Q(Q[12]) );
  FD_52 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n2), .Q(Q[13]) );
  FD_51 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n2), .Q(Q[14]) );
  FD_50 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n2), .Q(Q[15]) );
  FD_49 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n2), .Q(Q[16]) );
  FD_48 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n2), .Q(Q[17]) );
  FD_47 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n2), .Q(Q[18]) );
  FD_46 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n2), .Q(Q[19]) );
  FD_45 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n2), .Q(Q[20]) );
  FD_44 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n2), .Q(Q[21]) );
  FD_43 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n2), .Q(Q[22]) );
  FD_42 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n2), .Q(Q[23]) );
  FD_41 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n3), .Q(Q[24]) );
  FD_40 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n3), .Q(Q[25]) );
  FD_39 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n3), .Q(Q[26]) );
  FD_38 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n3), .Q(Q[27]) );
  FD_37 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n3), .Q(Q[28]) );
  FD_36 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n3), .Q(Q[29]) );
  FD_35 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n3), .Q(Q[30]) );
  FD_34 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n1) );
  BUF_X1 U2 ( .A(RESET), .Z(n2) );
  BUF_X1 U3 ( .A(RESET), .Z(n3) );
endmodule


module FD_33 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_32 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_31 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_30 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_29 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X2 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_28 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_27 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_26 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_25 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_24 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_23 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_22 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_21 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_20 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_19 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_18 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_17 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_16 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_15 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_14 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_13 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n1) );
endmodule


module FD_12 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_11 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_10 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_9 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_8 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(RESET), .ZN(n1) );
  AND2_X1 U4 ( .A1(D), .A2(n1), .ZN(N3) );
endmodule


module FD_7 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(D), .A2(n1), .ZN(N3) );
  INV_X1 U4 ( .A(RESET), .ZN(n1) );
endmodule


module FD_6 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_5 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X2 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(RESET), .ZN(n1) );
  AND2_X1 U4 ( .A1(D), .A2(n1), .ZN(N3) );
endmodule


module FD_4 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_3 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(RESET), .ZN(n1) );
  AND2_X1 U4 ( .A1(D), .A2(n1), .ZN(N3) );
endmodule


module FD_2 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_1 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n1;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(RESET), .ZN(N3) );
endmodule


module FD_GENERIC_NBIT33 ( D, CLK, RESET, Q );
  input [32:0] D;
  output [32:0] Q;
  input CLK, RESET;
  wire   n1, n2, n3;

  FD_33 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n1), .Q(Q[0]) );
  FD_32 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n1), .Q(Q[1]) );
  FD_31 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n1), .Q(Q[2]) );
  FD_30 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n1), .Q(Q[3]) );
  FD_29 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n1), .Q(Q[4]) );
  FD_28 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n1), .Q(Q[5]) );
  FD_27 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n1), .Q(Q[6]) );
  FD_26 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n1), .Q(Q[7]) );
  FD_25 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n1), .Q(Q[8]) );
  FD_24 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n1), .Q(Q[9]) );
  FD_23 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n1), .Q(Q[10]) );
  FD_22 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n1), .Q(Q[11]) );
  FD_21 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n2), .Q(Q[12]) );
  FD_20 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n2), .Q(Q[13]) );
  FD_19 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n2), .Q(Q[14]) );
  FD_18 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n2), .Q(Q[15]) );
  FD_17 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n2), .Q(Q[16]) );
  FD_16 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n2), .Q(Q[17]) );
  FD_15 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n2), .Q(Q[18]) );
  FD_14 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n2), .Q(Q[19]) );
  FD_13 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n2), .Q(Q[20]) );
  FD_12 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n2), .Q(Q[21]) );
  FD_11 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n2), .Q(Q[22]) );
  FD_10 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n2), .Q(Q[23]) );
  FD_9 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n2), .Q(Q[24]) );
  FD_8 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n3), .Q(Q[25]) );
  FD_7 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n3), .Q(Q[26]) );
  FD_6 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n3), .Q(Q[27]) );
  FD_5 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n3), .Q(Q[28]) );
  FD_4 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n3), .Q(Q[29]) );
  FD_3 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n3), .Q(Q[30]) );
  FD_2 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n3), .Q(Q[31]) );
  FD_1 FD_i_32 ( .D(D[32]), .CLK(CLK), .RESET(n3), .Q(Q[32]) );
  BUF_X1 U1 ( .A(RESET), .Z(n3) );
  BUF_X1 U2 ( .A(RESET), .Z(n1) );
  BUF_X1 U3 ( .A(RESET), .Z(n2) );
endmodule


module G_block_0 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1329, n1;
  assign G_OUT = net1329;

  AOI21_X1 U1 ( .B1(PG_IN_1), .B2(G_IN), .A(PG_IN_2), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net1329) );
endmodule


module G_block_9 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1440, n1, n2, n3;
  assign G_OUT = net1440;

  NOR2_X1 U1 ( .A1(PG_IN_1), .A2(PG_IN_2), .ZN(n3) );
  AOI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(net1440) );
  INV_X1 U3 ( .A(G_IN), .ZN(n1) );
  INV_X1 U4 ( .A(PG_IN_2), .ZN(n2) );
endmodule


module G_block_8 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(n2), .A2(n3), .ZN(G_OUT) );
  NAND2_X1 U2 ( .A1(G_IN), .A2(PG_IN_1), .ZN(n2) );
  INV_X1 U3 ( .A(PG_IN_2), .ZN(n3) );
endmodule


module G_block_7 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1603, n1;
  assign G_OUT = net1603;

  AOI21_X1 U1 ( .B1(G_IN), .B2(PG_IN_1), .A(PG_IN_2), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net1603) );
endmodule


module G_block_6 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_OUT) );
  AOI21_X1 U2 ( .B1(G_IN), .B2(PG_IN_1), .A(PG_IN_2), .ZN(n3) );
endmodule


module G_block_5 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1597, n1;
  assign G_OUT = net1597;

  INV_X1 U1 ( .A(n1), .ZN(net1597) );
  AOI21_X1 U2 ( .B1(G_IN), .B2(PG_IN_1), .A(PG_IN_2), .ZN(n1) );
endmodule


module G_block_4 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1615, n1;
  assign G_OUT = net1615;

  AOI21_X1 U1 ( .B1(G_IN), .B2(PG_IN_1), .A(PG_IN_2), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net1615) );
endmodule


module G_block_3 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1621, n1;
  assign G_OUT = net1621;

  OAI22_X1 U1 ( .A1(PG_IN_2), .A2(G_IN), .B1(PG_IN_1), .B2(PG_IN_2), .ZN(n1)
         );
  INV_X1 U2 ( .A(n1), .ZN(net1621) );
endmodule


module G_block_2 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   net1627, n1, n2;
  assign G_OUT = net1627;

  OR2_X1 U1 ( .A1(G_IN), .A2(PG_IN_2), .ZN(n1) );
  AND2_X2 U2 ( .A1(n1), .A2(n2), .ZN(net1627) );
  OR2_X1 U3 ( .A1(PG_IN_1), .A2(PG_IN_2), .ZN(n2) );
endmodule


module G_block_1 ( PG_IN_1, PG_IN_2, G_IN, G_OUT );
  input PG_IN_1, PG_IN_2, G_IN;
  output G_OUT;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_OUT) );
  AOI21_X1 U2 ( .B1(G_IN), .B2(PG_IN_1), .A(PG_IN_2), .ZN(n3) );
endmodule


module PG_block_0 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n1;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(PG_OUT_G) );
endmodule


module PG_block_26 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_25 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n1;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(PG_OUT_G) );
endmodule


module PG_block_24 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_23 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_22 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_21 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n1, n2, n3;

  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(PG_OUT_G) );
  INV_X1 U2 ( .A(PG_IN_first_G), .ZN(n1) );
  INV_X1 U3 ( .A(PG_IN_second_P), .ZN(n2) );
  INV_X1 U4 ( .A(PG_IN_second_G), .ZN(n3) );
  AND2_X1 U5 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_20 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_19 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_18 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  INV_X1 U2 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U3 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
endmodule


module PG_block_17 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_16 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_15 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_14 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_13 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_12 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n1;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(PG_OUT_G) );
endmodule


module PG_block_11 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n1, n2, n3;

  OAI21_X1 U1 ( .B1(n1), .B2(n2), .A(n3), .ZN(PG_OUT_G) );
  INV_X1 U2 ( .A(PG_IN_first_G), .ZN(n1) );
  INV_X1 U3 ( .A(PG_IN_second_P), .ZN(n2) );
  INV_X1 U4 ( .A(PG_IN_second_G), .ZN(n3) );
  AND2_X1 U5 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_10 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_9 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_8 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_7 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  INV_X1 U2 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U3 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
endmodule


module PG_block_6 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_5 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(PG_OUT_G) );
endmodule


module PG_block_4 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_3 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U2 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
  AND2_X1 U3 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
endmodule


module PG_block_2 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  INV_X1 U2 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U3 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
endmodule


module PG_block_1 ( PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, 
        PG_IN_second_G, PG_OUT_G, PG_OUT_PG );
  input PG_IN_first_P, PG_IN_second_P, PG_IN_first_G, PG_IN_second_G;
  output PG_OUT_G, PG_OUT_PG;
  wire   n3;

  AND2_X1 U1 ( .A1(PG_IN_second_P), .A2(PG_IN_first_P), .ZN(PG_OUT_PG) );
  INV_X1 U2 ( .A(n3), .ZN(PG_OUT_G) );
  AOI21_X1 U3 ( .B1(PG_IN_first_G), .B2(PG_IN_second_P), .A(PG_IN_second_G), 
        .ZN(n3) );
endmodule


module carry_generator_NBIT_GEN32_NBIT_Co8_N_ITERATION5 ( ADD_1, ADD_2, 
        Ci_carry_gen, Co );
  input [31:0] ADD_1;
  input [31:0] ADD_2;
  output [8:0] Co;
  input Ci_carry_gen;
  wire   Ci_carry_gen, n6, n7, n8, \G_matrix[15][15] , \G_matrix[15][14] ,
         \G_matrix[15][12] , \G_matrix[15][8] , \G_matrix[14][14] ,
         \G_matrix[13][13] , \G_matrix[13][12] , \G_matrix[12][12] ,
         \G_matrix[11][11] , \G_matrix[11][10] , \G_matrix[11][8] ,
         \G_matrix[10][10] , \G_matrix[9][9] , \G_matrix[9][8] ,
         \G_matrix[8][8] , \G_matrix[7][7] , \G_matrix[7][6] ,
         \G_matrix[7][4] , \G_matrix[6][6] , \G_matrix[5][5] ,
         \G_matrix[5][4] , \G_matrix[4][4] , \G_matrix[3][3] ,
         \G_matrix[3][2] , \G_matrix[2][2] , \G_matrix[2][0] ,
         \G_matrix[1][1] , \G_matrix[1][0] , \G_matrix[0][0] ,
         \G_matrix[31][31] , \G_matrix[31][30] , \G_matrix[31][28] ,
         \G_matrix[31][24] , \G_matrix[31][16] , \G_matrix[30][30] ,
         \G_matrix[29][29] , \G_matrix[29][28] , \G_matrix[28][28] ,
         \G_matrix[27][27] , \G_matrix[27][26] , \G_matrix[27][24] ,
         \G_matrix[27][16] , \G_matrix[26][26] , \G_matrix[25][25] ,
         \G_matrix[25][24] , \G_matrix[24][24] , \G_matrix[23][23] ,
         \G_matrix[23][22] , \G_matrix[23][20] , \G_matrix[23][16] ,
         \G_matrix[22][22] , \G_matrix[21][21] , \G_matrix[21][20] ,
         \G_matrix[20][20] , \G_matrix[19][19] , \G_matrix[19][18] ,
         \G_matrix[19][16] , \G_matrix[18][18] , \G_matrix[17][17] ,
         \G_matrix[17][16] , \G_matrix[16][16] , \PG_matrix[15][15] ,
         \PG_matrix[15][14] , \PG_matrix[15][12] , \PG_matrix[15][8] ,
         \PG_matrix[14][14] , \PG_matrix[13][13] , \PG_matrix[13][12] ,
         \PG_matrix[12][12] , \PG_matrix[11][11] , \PG_matrix[11][10] ,
         \PG_matrix[11][8] , \PG_matrix[10][10] , \PG_matrix[9][9] ,
         \PG_matrix[9][8] , \PG_matrix[8][8] , \PG_matrix[7][7] ,
         \PG_matrix[7][6] , \PG_matrix[7][4] , \PG_matrix[6][6] ,
         \PG_matrix[5][5] , \PG_matrix[5][4] , \PG_matrix[4][4] ,
         \PG_matrix[3][3] , \PG_matrix[3][2] , \PG_matrix[2][2] ,
         \PG_matrix[1][1] , \PG_matrix[0][0] , \PG_matrix[31][31] ,
         \PG_matrix[31][30] , \PG_matrix[31][28] , \PG_matrix[31][24] ,
         \PG_matrix[31][16] , \PG_matrix[30][30] , \PG_matrix[29][29] ,
         \PG_matrix[29][28] , \PG_matrix[28][28] , \PG_matrix[27][27] ,
         \PG_matrix[27][26] , \PG_matrix[27][24] , \PG_matrix[27][16] ,
         \PG_matrix[26][26] , \PG_matrix[25][25] , \PG_matrix[25][24] ,
         \PG_matrix[24][24] , \PG_matrix[23][23] , \PG_matrix[23][22] ,
         \PG_matrix[23][20] , \PG_matrix[23][16] , \PG_matrix[22][22] ,
         \PG_matrix[21][21] , \PG_matrix[21][20] , \PG_matrix[20][20] ,
         \PG_matrix[19][19] , \PG_matrix[19][18] , \PG_matrix[19][16] ,
         \PG_matrix[18][18] , \PG_matrix[17][17] , \PG_matrix[17][16] ,
         \PG_matrix[16][16] , net2479, net2480, n2, n4;
  assign Co[0] = Ci_carry_gen;

  XOR2_X1 U33 ( .A(ADD_2[9]), .B(ADD_1[9]), .Z(\PG_matrix[9][9] ) );
  XOR2_X1 U34 ( .A(ADD_2[8]), .B(ADD_1[8]), .Z(\PG_matrix[8][8] ) );
  XOR2_X1 U36 ( .A(ADD_2[6]), .B(ADD_1[6]), .Z(\PG_matrix[6][6] ) );
  XOR2_X1 U37 ( .A(ADD_2[5]), .B(ADD_1[5]), .Z(\PG_matrix[5][5] ) );
  XOR2_X1 U38 ( .A(ADD_2[4]), .B(ADD_1[4]), .Z(\PG_matrix[4][4] ) );
  XOR2_X1 U40 ( .A(ADD_2[31]), .B(ADD_1[31]), .Z(\PG_matrix[31][31] ) );
  XOR2_X1 U41 ( .A(ADD_2[30]), .B(ADD_1[30]), .Z(\PG_matrix[30][30] ) );
  XOR2_X1 U42 ( .A(ADD_2[2]), .B(ADD_1[2]), .Z(\PG_matrix[2][2] ) );
  XOR2_X1 U43 ( .A(ADD_2[29]), .B(ADD_1[29]), .Z(\PG_matrix[29][29] ) );
  XOR2_X1 U44 ( .A(ADD_2[28]), .B(ADD_1[28]), .Z(\PG_matrix[28][28] ) );
  XOR2_X1 U45 ( .A(ADD_2[27]), .B(ADD_1[27]), .Z(\PG_matrix[27][27] ) );
  XOR2_X1 U46 ( .A(ADD_2[26]), .B(ADD_1[26]), .Z(\PG_matrix[26][26] ) );
  XOR2_X1 U47 ( .A(ADD_2[25]), .B(ADD_1[25]), .Z(\PG_matrix[25][25] ) );
  XOR2_X1 U48 ( .A(ADD_2[24]), .B(ADD_1[24]), .Z(\PG_matrix[24][24] ) );
  XOR2_X1 U49 ( .A(ADD_2[23]), .B(ADD_1[23]), .Z(\PG_matrix[23][23] ) );
  XOR2_X1 U50 ( .A(ADD_2[22]), .B(ADD_1[22]), .Z(\PG_matrix[22][22] ) );
  XOR2_X1 U51 ( .A(ADD_2[21]), .B(ADD_1[21]), .Z(\PG_matrix[21][21] ) );
  XOR2_X1 U52 ( .A(ADD_2[20]), .B(ADD_1[20]), .Z(\PG_matrix[20][20] ) );
  XOR2_X1 U53 ( .A(ADD_2[1]), .B(ADD_1[1]), .Z(\PG_matrix[1][1] ) );
  XOR2_X1 U54 ( .A(ADD_2[19]), .B(ADD_1[19]), .Z(\PG_matrix[19][19] ) );
  XOR2_X1 U55 ( .A(ADD_2[18]), .B(ADD_1[18]), .Z(\PG_matrix[18][18] ) );
  XOR2_X1 U56 ( .A(ADD_2[17]), .B(ADD_1[17]), .Z(\PG_matrix[17][17] ) );
  XOR2_X1 U57 ( .A(ADD_2[16]), .B(ADD_1[16]), .Z(\PG_matrix[16][16] ) );
  XOR2_X1 U58 ( .A(ADD_2[15]), .B(ADD_1[15]), .Z(\PG_matrix[15][15] ) );
  XOR2_X1 U59 ( .A(ADD_2[14]), .B(ADD_1[14]), .Z(\PG_matrix[14][14] ) );
  XOR2_X1 U60 ( .A(ADD_2[13]), .B(ADD_1[13]), .Z(\PG_matrix[13][13] ) );
  XOR2_X1 U61 ( .A(ADD_2[12]), .B(ADD_1[12]), .Z(\PG_matrix[12][12] ) );
  XOR2_X1 U62 ( .A(ADD_2[11]), .B(ADD_1[11]), .Z(\PG_matrix[11][11] ) );
  XOR2_X1 U63 ( .A(ADD_2[10]), .B(ADD_1[10]), .Z(\PG_matrix[10][10] ) );
  G_block_0 G_block_0 ( .PG_IN_1(\PG_matrix[0][0] ), .PG_IN_2(\G_matrix[0][0] ), .G_IN(Ci_carry_gen), .G_OUT(\G_matrix[1][0] ) );
  G_block_9 G_block_2_0 ( .PG_IN_1(\PG_matrix[1][1] ), .PG_IN_2(
        \G_matrix[1][1] ), .G_IN(\G_matrix[1][0] ), .G_OUT(\G_matrix[2][0] )
         );
  G_block_8 G_block_3_0 ( .PG_IN_1(\PG_matrix[3][2] ), .PG_IN_2(
        \G_matrix[3][2] ), .G_IN(\G_matrix[2][0] ), .G_OUT(n8) );
  G_block_7 G_block_7_1 ( .PG_IN_1(\PG_matrix[7][4] ), .PG_IN_2(
        \G_matrix[7][4] ), .G_IN(n8), .G_OUT(n7) );
  G_block_6 G_block_cycle_2_1 ( .PG_IN_1(\PG_matrix[11][8] ), .PG_IN_2(
        \G_matrix[11][8] ), .G_IN(n4), .G_OUT(Co[3]) );
  G_block_5 G_block_cycle_2_2 ( .PG_IN_1(\PG_matrix[15][8] ), .PG_IN_2(
        \G_matrix[15][8] ), .G_IN(n7), .G_OUT(n6) );
  G_block_4 G_block_cycle_3_1 ( .PG_IN_1(\PG_matrix[19][16] ), .PG_IN_2(
        \G_matrix[19][16] ), .G_IN(n6), .G_OUT(Co[5]) );
  G_block_3 G_block_cycle_3_2 ( .PG_IN_1(\PG_matrix[23][16] ), .PG_IN_2(n2), 
        .G_IN(n6), .G_OUT(Co[6]) );
  G_block_2 G_block_cycle_3_3 ( .PG_IN_1(\PG_matrix[27][16] ), .PG_IN_2(
        \G_matrix[27][16] ), .G_IN(n6), .G_OUT(Co[7]) );
  G_block_1 G_block_cycle_3_4 ( .PG_IN_1(\PG_matrix[31][16] ), .PG_IN_2(
        \G_matrix[31][16] ), .G_IN(Co[4]), .G_OUT(Co[8]) );
  PG_block_0 pre_generation_0_1 ( .PG_IN_first_P(\PG_matrix[2][2] ), 
        .PG_IN_second_P(\PG_matrix[3][3] ), .PG_IN_first_G(\G_matrix[2][2] ), 
        .PG_IN_second_G(\G_matrix[3][3] ), .PG_OUT_G(\G_matrix[3][2] ), 
        .PG_OUT_PG(\PG_matrix[3][2] ) );
  PG_block_26 pre_generation_0_2 ( .PG_IN_first_P(\PG_matrix[4][4] ), 
        .PG_IN_second_P(\PG_matrix[5][5] ), .PG_IN_first_G(\G_matrix[4][4] ), 
        .PG_IN_second_G(\G_matrix[5][5] ), .PG_OUT_G(\G_matrix[5][4] ), 
        .PG_OUT_PG(\PG_matrix[5][4] ) );
  PG_block_25 pre_generation_0_3 ( .PG_IN_first_P(\PG_matrix[6][6] ), 
        .PG_IN_second_P(\PG_matrix[7][7] ), .PG_IN_first_G(\G_matrix[6][6] ), 
        .PG_IN_second_G(\G_matrix[7][7] ), .PG_OUT_G(\G_matrix[7][6] ), 
        .PG_OUT_PG(\PG_matrix[7][6] ) );
  PG_block_24 pre_generation_0_4 ( .PG_IN_first_P(\PG_matrix[8][8] ), 
        .PG_IN_second_P(\PG_matrix[9][9] ), .PG_IN_first_G(\G_matrix[8][8] ), 
        .PG_IN_second_G(\G_matrix[9][9] ), .PG_OUT_G(\G_matrix[9][8] ), 
        .PG_OUT_PG(\PG_matrix[9][8] ) );
  PG_block_23 pre_generation_0_5 ( .PG_IN_first_P(\PG_matrix[10][10] ), 
        .PG_IN_second_P(\PG_matrix[11][11] ), .PG_IN_first_G(
        \G_matrix[10][10] ), .PG_IN_second_G(\G_matrix[11][11] ), .PG_OUT_G(
        \G_matrix[11][10] ), .PG_OUT_PG(\PG_matrix[11][10] ) );
  PG_block_22 pre_generation_0_6 ( .PG_IN_first_P(\PG_matrix[12][12] ), 
        .PG_IN_second_P(\PG_matrix[13][13] ), .PG_IN_first_G(
        \G_matrix[12][12] ), .PG_IN_second_G(\G_matrix[13][13] ), .PG_OUT_G(
        \G_matrix[13][12] ), .PG_OUT_PG(\PG_matrix[13][12] ) );
  PG_block_21 pre_generation_0_7 ( .PG_IN_first_P(\PG_matrix[14][14] ), 
        .PG_IN_second_P(\PG_matrix[15][15] ), .PG_IN_first_G(
        \G_matrix[14][14] ), .PG_IN_second_G(\G_matrix[15][15] ), .PG_OUT_G(
        \G_matrix[15][14] ), .PG_OUT_PG(\PG_matrix[15][14] ) );
  PG_block_20 pre_generation_0_8 ( .PG_IN_first_P(\PG_matrix[16][16] ), 
        .PG_IN_second_P(\PG_matrix[17][17] ), .PG_IN_first_G(
        \G_matrix[16][16] ), .PG_IN_second_G(\G_matrix[17][17] ), .PG_OUT_G(
        \G_matrix[17][16] ), .PG_OUT_PG(\PG_matrix[17][16] ) );
  PG_block_19 pre_generation_0_9 ( .PG_IN_first_P(\PG_matrix[18][18] ), 
        .PG_IN_second_P(\PG_matrix[19][19] ), .PG_IN_first_G(
        \G_matrix[18][18] ), .PG_IN_second_G(\G_matrix[19][19] ), .PG_OUT_G(
        \G_matrix[19][18] ), .PG_OUT_PG(\PG_matrix[19][18] ) );
  PG_block_18 pre_generation_0_10 ( .PG_IN_first_P(\PG_matrix[20][20] ), 
        .PG_IN_second_P(\PG_matrix[21][21] ), .PG_IN_first_G(
        \G_matrix[20][20] ), .PG_IN_second_G(\G_matrix[21][21] ), .PG_OUT_G(
        \G_matrix[21][20] ), .PG_OUT_PG(\PG_matrix[21][20] ) );
  PG_block_17 pre_generation_0_11 ( .PG_IN_first_P(\PG_matrix[22][22] ), 
        .PG_IN_second_P(\PG_matrix[23][23] ), .PG_IN_first_G(
        \G_matrix[22][22] ), .PG_IN_second_G(\G_matrix[23][23] ), .PG_OUT_G(
        \G_matrix[23][22] ), .PG_OUT_PG(\PG_matrix[23][22] ) );
  PG_block_16 pre_generation_0_12 ( .PG_IN_first_P(\PG_matrix[24][24] ), 
        .PG_IN_second_P(\PG_matrix[25][25] ), .PG_IN_first_G(
        \G_matrix[24][24] ), .PG_IN_second_G(\G_matrix[25][25] ), .PG_OUT_G(
        \G_matrix[25][24] ), .PG_OUT_PG(\PG_matrix[25][24] ) );
  PG_block_15 pre_generation_0_13 ( .PG_IN_first_P(\PG_matrix[26][26] ), 
        .PG_IN_second_P(\PG_matrix[27][27] ), .PG_IN_first_G(
        \G_matrix[26][26] ), .PG_IN_second_G(\G_matrix[27][27] ), .PG_OUT_G(
        \G_matrix[27][26] ), .PG_OUT_PG(\PG_matrix[27][26] ) );
  PG_block_14 pre_generation_0_14 ( .PG_IN_first_P(\PG_matrix[28][28] ), 
        .PG_IN_second_P(\PG_matrix[29][29] ), .PG_IN_first_G(
        \G_matrix[28][28] ), .PG_IN_second_G(\G_matrix[29][29] ), .PG_OUT_G(
        \G_matrix[29][28] ), .PG_OUT_PG(\PG_matrix[29][28] ) );
  PG_block_13 pre_generation_0_15 ( .PG_IN_first_P(\PG_matrix[30][30] ), 
        .PG_IN_second_P(\PG_matrix[31][31] ), .PG_IN_first_G(
        \G_matrix[30][30] ), .PG_IN_second_G(\G_matrix[31][31] ), .PG_OUT_G(
        \G_matrix[31][30] ), .PG_OUT_PG(\PG_matrix[31][30] ) );
  PG_block_12 pre_generation_1_0 ( .PG_IN_first_P(\PG_matrix[5][4] ), 
        .PG_IN_second_P(\PG_matrix[7][6] ), .PG_IN_first_G(\G_matrix[5][4] ), 
        .PG_IN_second_G(\G_matrix[7][6] ), .PG_OUT_G(\G_matrix[7][4] ), 
        .PG_OUT_PG(\PG_matrix[7][4] ) );
  PG_block_11 pre_generation_1_1 ( .PG_IN_first_P(\PG_matrix[9][8] ), 
        .PG_IN_second_P(\PG_matrix[11][10] ), .PG_IN_first_G(\G_matrix[9][8] ), 
        .PG_IN_second_G(\G_matrix[11][10] ), .PG_OUT_G(\G_matrix[11][8] ), 
        .PG_OUT_PG(\PG_matrix[11][8] ) );
  PG_block_10 pre_generation_1_2 ( .PG_IN_first_P(\PG_matrix[13][12] ), 
        .PG_IN_second_P(\PG_matrix[15][14] ), .PG_IN_first_G(
        \G_matrix[13][12] ), .PG_IN_second_G(\G_matrix[15][14] ), .PG_OUT_G(
        \G_matrix[15][12] ), .PG_OUT_PG(\PG_matrix[15][12] ) );
  PG_block_9 pre_generation_1_3 ( .PG_IN_first_P(\PG_matrix[17][16] ), 
        .PG_IN_second_P(\PG_matrix[19][18] ), .PG_IN_first_G(
        \G_matrix[17][16] ), .PG_IN_second_G(\G_matrix[19][18] ), .PG_OUT_G(
        \G_matrix[19][16] ), .PG_OUT_PG(\PG_matrix[19][16] ) );
  PG_block_8 pre_generation_1_4 ( .PG_IN_first_P(\PG_matrix[21][20] ), 
        .PG_IN_second_P(\PG_matrix[23][22] ), .PG_IN_first_G(
        \G_matrix[21][20] ), .PG_IN_second_G(\G_matrix[23][22] ), .PG_OUT_G(
        \G_matrix[23][20] ), .PG_OUT_PG(\PG_matrix[23][20] ) );
  PG_block_7 pre_generation_1_5 ( .PG_IN_first_P(\PG_matrix[25][24] ), 
        .PG_IN_second_P(\PG_matrix[27][26] ), .PG_IN_first_G(
        \G_matrix[25][24] ), .PG_IN_second_G(\G_matrix[27][26] ), .PG_OUT_G(
        \G_matrix[27][24] ), .PG_OUT_PG(\PG_matrix[27][24] ) );
  PG_block_6 pre_generation_1_6 ( .PG_IN_first_P(\PG_matrix[29][28] ), 
        .PG_IN_second_P(\PG_matrix[31][30] ), .PG_IN_first_G(
        \G_matrix[29][28] ), .PG_IN_second_G(\G_matrix[31][30] ), .PG_OUT_G(
        \G_matrix[31][28] ), .PG_OUT_PG(\PG_matrix[31][28] ) );
  PG_block_5 gen_2_0_0 ( .PG_IN_first_P(\PG_matrix[11][8] ), .PG_IN_second_P(
        \PG_matrix[15][12] ), .PG_IN_first_G(\G_matrix[11][8] ), 
        .PG_IN_second_G(\G_matrix[15][12] ), .PG_OUT_G(\G_matrix[15][8] ), 
        .PG_OUT_PG(\PG_matrix[15][8] ) );
  PG_block_4 gen_2_0_1 ( .PG_IN_first_P(\PG_matrix[19][16] ), .PG_IN_second_P(
        \PG_matrix[23][20] ), .PG_IN_first_G(\G_matrix[19][16] ), 
        .PG_IN_second_G(\G_matrix[23][20] ), .PG_OUT_G(\G_matrix[23][16] ), 
        .PG_OUT_PG(\PG_matrix[23][16] ) );
  PG_block_3 gen_2_0_2 ( .PG_IN_first_P(\PG_matrix[27][24] ), .PG_IN_second_P(
        \PG_matrix[31][28] ), .PG_IN_first_G(\G_matrix[27][24] ), 
        .PG_IN_second_G(\G_matrix[31][28] ), .PG_OUT_G(\G_matrix[31][24] ), 
        .PG_OUT_PG(\PG_matrix[31][24] ) );
  PG_block_2 PG_block_cycle_1_1_1 ( .PG_IN_first_P(\PG_matrix[23][16] ), 
        .PG_IN_second_P(\PG_matrix[27][24] ), .PG_IN_first_G(
        \G_matrix[23][16] ), .PG_IN_second_G(\G_matrix[27][24] ), .PG_OUT_G(
        \G_matrix[27][16] ), .PG_OUT_PG(\PG_matrix[27][16] ) );
  PG_block_1 PG_block_cycle_1_1_2 ( .PG_IN_first_P(\PG_matrix[23][16] ), 
        .PG_IN_second_P(\PG_matrix[31][24] ), .PG_IN_first_G(n2), 
        .PG_IN_second_G(\G_matrix[31][24] ), .PG_OUT_G(\G_matrix[31][16] ), 
        .PG_OUT_PG(\PG_matrix[31][16] ) );
  CLKBUF_X1 U1 ( .A(n6), .Z(Co[4]) );
  BUF_X1 U2 ( .A(n4), .Z(Co[2]) );
  CLKBUF_X1 U3 ( .A(n7), .Z(n4) );
  CLKBUF_X1 U4 ( .A(\G_matrix[23][16] ), .Z(n2) );
  XOR2_X1 U5 ( .A(ADD_2[0]), .B(ADD_1[0]), .Z(\PG_matrix[0][0] ) );
  INV_X1 U6 ( .A(ADD_2[0]), .ZN(net2480) );
  INV_X1 U7 ( .A(ADD_1[0]), .ZN(net2479) );
  AND2_X1 U8 ( .A1(ADD_2[2]), .A2(ADD_1[2]), .ZN(\G_matrix[2][2] ) );
  AND2_X1 U9 ( .A1(ADD_2[3]), .A2(ADD_1[3]), .ZN(\G_matrix[3][3] ) );
  AND2_X1 U10 ( .A1(ADD_2[18]), .A2(ADD_1[18]), .ZN(\G_matrix[18][18] ) );
  AND2_X1 U11 ( .A1(ADD_2[19]), .A2(ADD_1[19]), .ZN(\G_matrix[19][19] ) );
  AND2_X1 U12 ( .A1(ADD_2[16]), .A2(ADD_1[16]), .ZN(\G_matrix[16][16] ) );
  AND2_X1 U13 ( .A1(ADD_2[17]), .A2(ADD_1[17]), .ZN(\G_matrix[17][17] ) );
  AND2_X1 U14 ( .A1(ADD_2[10]), .A2(ADD_1[10]), .ZN(\G_matrix[10][10] ) );
  AND2_X1 U15 ( .A1(ADD_2[11]), .A2(ADD_1[11]), .ZN(\G_matrix[11][11] ) );
  AND2_X1 U16 ( .A1(ADD_2[8]), .A2(ADD_1[8]), .ZN(\G_matrix[8][8] ) );
  AND2_X1 U17 ( .A1(ADD_2[9]), .A2(ADD_1[9]), .ZN(\G_matrix[9][9] ) );
  AND2_X1 U18 ( .A1(ADD_2[12]), .A2(ADD_1[12]), .ZN(\G_matrix[12][12] ) );
  AND2_X1 U19 ( .A1(ADD_2[13]), .A2(ADD_1[13]), .ZN(\G_matrix[13][13] ) );
  AND2_X1 U20 ( .A1(ADD_2[22]), .A2(ADD_1[22]), .ZN(\G_matrix[22][22] ) );
  AND2_X1 U21 ( .A1(ADD_2[23]), .A2(ADD_1[23]), .ZN(\G_matrix[23][23] ) );
  AND2_X1 U22 ( .A1(ADD_2[4]), .A2(ADD_1[4]), .ZN(\G_matrix[4][4] ) );
  AND2_X1 U23 ( .A1(ADD_2[5]), .A2(ADD_1[5]), .ZN(\G_matrix[5][5] ) );
  AND2_X1 U24 ( .A1(ADD_2[26]), .A2(ADD_1[26]), .ZN(\G_matrix[26][26] ) );
  AND2_X1 U25 ( .A1(ADD_2[27]), .A2(ADD_1[27]), .ZN(\G_matrix[27][27] ) );
  AND2_X1 U26 ( .A1(ADD_2[24]), .A2(ADD_1[24]), .ZN(\G_matrix[24][24] ) );
  AND2_X1 U27 ( .A1(ADD_2[25]), .A2(ADD_1[25]), .ZN(\G_matrix[25][25] ) );
  AND2_X1 U28 ( .A1(ADD_2[30]), .A2(ADD_1[30]), .ZN(\G_matrix[30][30] ) );
  AND2_X1 U29 ( .A1(ADD_2[31]), .A2(ADD_1[31]), .ZN(\G_matrix[31][31] ) );
  AND2_X1 U30 ( .A1(ADD_2[29]), .A2(ADD_1[29]), .ZN(\G_matrix[29][29] ) );
  AND2_X1 U31 ( .A1(ADD_2[28]), .A2(ADD_1[28]), .ZN(\G_matrix[28][28] ) );
  AND2_X1 U32 ( .A1(ADD_2[14]), .A2(ADD_1[14]), .ZN(\G_matrix[14][14] ) );
  AND2_X1 U35 ( .A1(ADD_2[15]), .A2(ADD_1[15]), .ZN(\G_matrix[15][15] ) );
  AND2_X1 U39 ( .A1(ADD_2[1]), .A2(ADD_1[1]), .ZN(\G_matrix[1][1] ) );
  AND2_X1 U64 ( .A1(ADD_2[20]), .A2(ADD_1[20]), .ZN(\G_matrix[20][20] ) );
  AND2_X1 U65 ( .A1(ADD_2[21]), .A2(ADD_1[21]), .ZN(\G_matrix[21][21] ) );
  AND2_X1 U66 ( .A1(ADD_2[6]), .A2(ADD_1[6]), .ZN(\G_matrix[6][6] ) );
  AND2_X1 U67 ( .A1(ADD_2[7]), .A2(ADD_1[7]), .ZN(\G_matrix[7][7] ) );
  CLKBUF_X1 U68 ( .A(n8), .Z(Co[1]) );
  XOR2_X1 U69 ( .A(ADD_2[7]), .B(ADD_1[7]), .Z(\PG_matrix[7][7] ) );
  XOR2_X1 U70 ( .A(ADD_2[3]), .B(ADD_1[3]), .Z(\PG_matrix[3][3] ) );
  NOR2_X1 U71 ( .A1(net2479), .A2(net2480), .ZN(\G_matrix[0][0] ) );
endmodule


module RCA_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(Ci), .B(B[0]), .CI(A[0]), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(Ci), .B(B[0]), .CI(A[0]), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n5;

  INV_X1 U1 ( .A(n9), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n6), .ZN(Y[3]) );
  INV_X1 U3 ( .A(n7), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n5), .ZN(n6) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n5), .ZN(n7) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n5), .ZN(n8) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n5), .ZN(n9) );
  INV_X1 U9 ( .A(SEL), .ZN(n5) );
endmodule


module carry_select_block_NBIT4_0 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_0 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_15 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_0 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n5, n10, n11, n12, n13;

  INV_X1 U1 ( .A(n10), .ZN(Y[0]) );
  INV_X1 U2 ( .A(n11), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n12), .ZN(Y[2]) );
  INV_X1 U4 ( .A(n13), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n13) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n5), .ZN(n12) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n5), .ZN(n11) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n5), .ZN(n10) );
  INV_X1 U9 ( .A(SEL), .ZN(n5) );
endmodule


module carry_select_block_NBIT4_7 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_14 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_13 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_7 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n10, n11, n12, n13, n14;

  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  INV_X1 U2 ( .A(n11), .ZN(Y[0]) );
  INV_X1 U3 ( .A(n12), .ZN(Y[1]) );
  INV_X1 U4 ( .A(n13), .ZN(Y[2]) );
  INV_X1 U5 ( .A(n14), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(n1), .A2(A[3]), .B1(B[3]), .B2(n10), .ZN(n14) );
  AOI22_X1 U7 ( .A1(n1), .A2(A[2]), .B1(B[2]), .B2(n10), .ZN(n13) );
  AOI22_X1 U8 ( .A1(n1), .A2(A[1]), .B1(B[1]), .B2(n10), .ZN(n12) );
  AOI22_X1 U9 ( .A1(n1), .A2(A[0]), .B1(B[0]), .B2(n10), .ZN(n11) );
  INV_X1 U10 ( .A(SEL), .ZN(n10) );
endmodule


module carry_select_block_NBIT4_6 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_12 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_11 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_6 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n11, n12, n13, n14, n15;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  INV_X1 U3 ( .A(SEL), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(Y[0]) );
  AOI22_X1 U5 ( .A1(n1), .A2(A[0]), .B1(n11), .B2(B[0]), .ZN(n12) );
  INV_X1 U6 ( .A(n13), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(n2), .A2(A[1]), .B1(n11), .B2(B[1]), .ZN(n13) );
  INV_X1 U8 ( .A(n15), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(n1), .A2(A[3]), .B1(n11), .B2(B[3]), .ZN(n15) );
  INV_X1 U10 ( .A(n14), .ZN(Y[2]) );
  AOI22_X1 U11 ( .A1(n2), .A2(A[2]), .B1(n11), .B2(B[2]), .ZN(n14) );
endmodule


module carry_select_block_NBIT4_5 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_10 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_9 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_5 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n12, n13, n14, n15;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  INV_X1 U3 ( .A(SEL), .ZN(n3) );
  INV_X1 U4 ( .A(n12), .ZN(Y[0]) );
  INV_X1 U5 ( .A(n13), .ZN(Y[1]) );
  INV_X1 U6 ( .A(n14), .ZN(Y[2]) );
  INV_X1 U7 ( .A(n15), .ZN(Y[3]) );
  AOI22_X1 U8 ( .A1(n2), .A2(A[3]), .B1(n3), .B2(B[3]), .ZN(n15) );
  AOI22_X1 U9 ( .A1(n2), .A2(A[2]), .B1(n3), .B2(B[2]), .ZN(n14) );
  AOI22_X1 U10 ( .A1(n1), .A2(A[1]), .B1(n3), .B2(B[1]), .ZN(n13) );
  AOI22_X1 U11 ( .A1(n1), .A2(A[0]), .B1(n3), .B2(B[0]), .ZN(n12) );
endmodule


module carry_select_block_NBIT4_4 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_8 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_7 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_4 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n5, n6, n8, n9, n11, n13, n14, n15, n16, n17;

  CLKBUF_X1 U1 ( .A(SEL), .Z(n17) );
  BUF_X1 U2 ( .A(SEL), .Z(n15) );
  BUF_X1 U3 ( .A(SEL), .Z(n1) );
  NAND2_X1 U4 ( .A1(n1), .A2(A[3]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n16), .A2(B[3]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(n3), .A2(n2), .ZN(Y[3]) );
  NAND2_X1 U7 ( .A1(n15), .A2(A[2]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(n16), .A2(B[2]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(n6), .A2(n5), .ZN(Y[2]) );
  NAND2_X1 U10 ( .A1(n1), .A2(A[1]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(n16), .A2(B[1]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(n9), .A2(n8), .ZN(Y[1]) );
  INV_X1 U13 ( .A(A[0]), .ZN(n13) );
  INV_X1 U14 ( .A(n17), .ZN(n11) );
  INV_X1 U15 ( .A(B[0]), .ZN(n14) );
  OAI22_X1 U16 ( .A1(n11), .A2(n13), .B1(n15), .B2(n14), .ZN(Y[0]) );
  INV_X1 U17 ( .A(SEL), .ZN(n16) );
endmodule


module carry_select_block_NBIT4_3 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_6 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_5 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_3 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   net1475, net2526, net2525, net2524, n2, n3, n5;
  assign Y[2] = net1475;
  assign Y[0] = net2524;

  MUX2_X1 U1 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
  NAND2_X1 U2 ( .A1(SEL), .A2(A[3]), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n5), .A2(B[3]), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Y[3]) );
  INV_X1 U5 ( .A(SEL), .ZN(n5) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(net1475) );
  OAI22_X1 U7 ( .A1(n5), .A2(net2525), .B1(SEL), .B2(net2526), .ZN(net2524) );
  INV_X1 U8 ( .A(B[0]), .ZN(net2526) );
  INV_X1 U9 ( .A(A[0]), .ZN(net2525) );
endmodule


module carry_select_block_NBIT4_2 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_4 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_3 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_2 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module RCA_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \r56/carry[3] , \r56/carry[2] , \r56/carry[1] ;

  FA_X1 \r56/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(\r56/carry[1] ), .S(S[0]) );
  FA_X1 \r56/U1_1  ( .A(A[1]), .B(B[1]), .CI(\r56/carry[1] ), .CO(
        \r56/carry[2] ), .S(S[1]) );
  FA_X1 \r56/U1_2  ( .A(A[2]), .B(B[2]), .CI(\r56/carry[2] ), .CO(
        \r56/carry[3] ), .S(S[2]) );
  FA_X1 \r56/U1_3  ( .A(A[3]), .B(B[3]), .CI(\r56/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   net1470, net2871, n1, n3;
  assign Y[2] = net1470;
  assign Y[0] = net2871;

  OAI21_X1 U1 ( .B1(SEL), .B2(n1), .A(n3), .ZN(Y[1]) );
  INV_X1 U2 ( .A(B[1]), .ZN(n1) );
  MUX2_X1 U3 ( .A(B[3]), .B(A[3]), .S(SEL), .Z(Y[3]) );
  NAND2_X1 U4 ( .A1(SEL), .A2(A[1]), .ZN(n3) );
  MUX2_X1 U5 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(net2871) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(net1470) );
endmodule


module carry_select_block_NBIT4_1 ( INPUT_1, INPUT_2, Ci_sel, SUM );
  input [3:0] INPUT_1;
  input [3:0] INPUT_2;
  output [3:0] SUM;
  input Ci_sel;

  wire   [3:0] SUM_0;
  wire   [3:0] SUM_1;

  RCA_NBIT4_2 ADDER0 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b0), .S(SUM_0) );
  RCA_NBIT4_1 ADDER1 ( .A(INPUT_1), .B(INPUT_2), .Ci(1'b1), .S(SUM_1) );
  MUX21_GENERIC_NBIT4_1 MUX ( .A(SUM_1), .B(SUM_0), .SEL(Ci_sel), .Y(SUM) );
endmodule


module sum_generator_NBIT_GEN32_NBIT_GEN_BLOCK8 ( ADD_1, ADD_2, Ci, SUM );
  input [31:0] ADD_1;
  input [31:0] ADD_2;
  input [7:0] Ci;
  output [31:0] SUM;


  carry_select_block_NBIT4_0 sum_gen_1 ( .INPUT_1(ADD_1[3:0]), .INPUT_2(
        ADD_2[3:0]), .Ci_sel(Ci[0]), .SUM(SUM[3:0]) );
  carry_select_block_NBIT4_7 sum_gen_2 ( .INPUT_1(ADD_1[7:4]), .INPUT_2(
        ADD_2[7:4]), .Ci_sel(Ci[1]), .SUM(SUM[7:4]) );
  carry_select_block_NBIT4_6 sum_gen_3 ( .INPUT_1(ADD_1[11:8]), .INPUT_2(
        ADD_2[11:8]), .Ci_sel(Ci[2]), .SUM(SUM[11:8]) );
  carry_select_block_NBIT4_5 sum_gen_4 ( .INPUT_1(ADD_1[15:12]), .INPUT_2(
        ADD_2[15:12]), .Ci_sel(Ci[3]), .SUM(SUM[15:12]) );
  carry_select_block_NBIT4_4 sum_gen_5 ( .INPUT_1(ADD_1[19:16]), .INPUT_2(
        ADD_2[19:16]), .Ci_sel(Ci[4]), .SUM(SUM[19:16]) );
  carry_select_block_NBIT4_3 sum_gen_6 ( .INPUT_1(ADD_1[23:20]), .INPUT_2(
        ADD_2[23:20]), .Ci_sel(Ci[5]), .SUM(SUM[23:20]) );
  carry_select_block_NBIT4_2 sum_gen_7 ( .INPUT_1(ADD_1[27:24]), .INPUT_2(
        ADD_2[27:24]), .Ci_sel(Ci[6]), .SUM(SUM[27:24]) );
  carry_select_block_NBIT4_1 sum_gen_8 ( .INPUT_1(ADD_1[31:28]), .INPUT_2(
        ADD_2[31:28]), .Ci_sel(Ci[7]), .SUM(SUM[31:28]) );
endmodule


module P4_adder_NBIT32 ( INPUT_1, INPUT_2, C_in, SUM, C_out, reset, Clk );
  input [31:0] INPUT_1;
  input [31:0] INPUT_2;
  output [32:0] SUM;
  input C_in, reset, Clk;
  output C_out;
  wire   n1, n2;
  wire   [31:0] in_1;
  wire   [31:0] in_2;
  wire   [7:0] Carry_from_carry_gen;
  wire   [32:1] p4_sum_and_cout;

  FD_GENERIC_NBIT32_0 reg_1 ( .D(INPUT_1), .CLK(Clk), .RESET(reset), .Q(in_1)
         );
  FD_GENERIC_NBIT32_1 reg_2 ( .D(INPUT_2), .CLK(Clk), .RESET(reset), .Q(in_2)
         );
  FD_GENERIC_NBIT33 reg_out ( .D({p4_sum_and_cout, C_out}), .CLK(Clk), .RESET(
        reset), .Q(SUM) );
  carry_generator_NBIT_GEN32_NBIT_Co8_N_ITERATION5 Carry_gen ( .ADD_1(in_1), 
        .ADD_2(in_2), .Ci_carry_gen(C_in), .Co({C_out, Carry_from_carry_gen})
         );
  sum_generator_NBIT_GEN32_NBIT_GEN_BLOCK8 Sum_gen ( .ADD_1({in_1[31:1], n2}), 
        .ADD_2({in_2[31:1], n1}), .Ci(Carry_from_carry_gen), .SUM(
        p4_sum_and_cout) );
  BUF_X1 U1 ( .A(in_2[0]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(in_1[0]), .Z(n2) );
endmodule

