
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_NBIT32_NADDRESS5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_NBIT32_NADDRESS5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_NBIT32_NADDRESS5.all;

entity register_file_NBIT32_NADDRESS5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT32_NADDRESS5;

architecture SYN_A of register_file_NBIT32_NADDRESS5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, 
      n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
      n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, 
      n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
      n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
      n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, 
      n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
      n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
      n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
      n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, 
      n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, 
      n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
      n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, 
      n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, 
      n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
      n2359, n2360, n2361, n2362, n2363, n12826, n12827, n12828, n12829, n12830
      , n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
      n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, 
      n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, 
      n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, 
      n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, 
      n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, 
      n12981, n12982, n12983, n12984, n12985, n13082, n13083, n13084, n13085, 
      n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, 
      n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, 
      n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, 
      n13113, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, 
      n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, 
      n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, 
      n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, 
      n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, 
      n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, 
      n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, 
      n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, 
      n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, 
      n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, 
      n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, 
      n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, 
      n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, 
      n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, 
      n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, 
      n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, 
      n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, 
      n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, 
      n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, 
      n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, 
      n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, 
      n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, 
      n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, 
      n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, 
      n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, 
      n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, 
      n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, 
      n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, 
      n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, 
      n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, 
      n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, 
      n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, 
      n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, 
      n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, 
      n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, 
      n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, 
      n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, 
      n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, 
      n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, 
      n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, 
      n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, 
      n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, 
      n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, 
      n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, 
      n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, 
      n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, 
      n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, 
      n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, 
      n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, 
      n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, 
      n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, 
      n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, 
      n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, 
      n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, 
      n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, 
      n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, 
      n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, 
      n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, 
      n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, 
      n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, 
      n13749, n13750, n13751, n13752, n13753, n14442, n14443, n14444, n14445, 
      n14446, n14447, n14450, n14451, n14452, n14453, n14454, n14457, n14458, 
      n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, 
      n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, 
      n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, 
      n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, 
      n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, 
      n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, 
      n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, 
      n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
      n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
      n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, 
      n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, 
      n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, 
      n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, 
      n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, 
      n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, 
      n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, 
      n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, 
      n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, 
      n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, 
      n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, 
      n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, 
      n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, 
      n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, 
      n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, 
      n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, 
      n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, 
      n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, 
      n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, 
      n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, 
      n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, 
      n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, 
      n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, 
      n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, 
      n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, 
      n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, 
      n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, 
      n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, 
      n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, 
      n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, 
      n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, 
      n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, 
      n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, 
      n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, 
      n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, 
      n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, 
      n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, 
      n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, 
      n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, 
      n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, 
      n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, 
      n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, 
      n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, 
      n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, 
      n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, 
      n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, 
      n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, 
      n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, 
      n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, 
      n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, 
      n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, 
      n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, 
      n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, 
      n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, 
      n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, 
      n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, 
      n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
      n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, 
      n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, 
      n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, 
      n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, 
      n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, 
      n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, 
      n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, 
      n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, 
      n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, 
      n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, 
      n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, 
      n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, 
      n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, 
      n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, 
      n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, 
      n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15226, 
      n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, 
      n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, 
      n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, 
      n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, 
      n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, 
      n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, 
      n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, 
      n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, 
      n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, 
      n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, 
      n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, 
      n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, 
      n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, 
      n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, 
      n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, 
      n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, 
      n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, 
      n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, 
      n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, 
      n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, 
      n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, 
      n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, 
      n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, 
      n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, 
      n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, 
      n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, 
      n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, 
      n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, 
      n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, 
      n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, 
      n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, 
      n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, 
      n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, 
      n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, 
      n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, 
      n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, 
      n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, 
      n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, 
      n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, 
      n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, 
      n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, 
      n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, 
      n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, 
      n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, 
      n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, 
      n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, 
      n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, 
      n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, 
      n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, 
      n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, 
      n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, 
      n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, 
      n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, 
      n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, 
      n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, 
      n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, 
      n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, 
      n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, 
      n15794, n15795, n15797, n15798, n15799, n15800, n15801, n15802, n15803, 
      n15804, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, 
      n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, 
      n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, 
      n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
      n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, 
      n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
      n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, 
      n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, 
      n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, 
      n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, 
      n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, 
      n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, 
      n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, 
      n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, 
      n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, 
      n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, 
      n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, 
      n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, 
      n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, 
      n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, 
      n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, 
      n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, 
      n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, 
      n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, 
      n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, 
      n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, 
      n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, 
      n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, 
      n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, 
      n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, 
      n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, 
      n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, 
      n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, 
      n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, 
      n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, 
      n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, 
      n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, 
      n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, 
      n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, 
      n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, 
      n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, 
      n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, 
      n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, 
      n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, 
      n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, 
      n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, 
      n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, 
      n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, 
      n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, 
      n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, 
      n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, 
      n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, 
      n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, 
      n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, 
      n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, 
      n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, 
      n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, 
      n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, 
      n16337, n16338, n16339, n16340, n16341, n16366, n16367, n16368, n16369, 
      n16370, n16371, n16372, n16373, n16382, n16383, n16384, n16385, n16386, 
      n16387, n16388, n16389, n16414, n16415, n16416, n16417, n16418, n16419, 
      n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, 
      n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, 
      n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, 
      n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, 
      n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, 
      n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, 
      n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, 
      n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, 
      n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, 
      n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, 
      n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, 
      n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16675, n16676, n16677, n16702, n16703, n16704, 
      n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, 
      n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, 
      n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, 
      n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, 
      n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, 
      n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, 
      n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, 
      n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, 
      n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, 
      n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, 
      n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, 
      n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, 
      n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, 
      n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, 
      n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, 
      n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, 
      n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, 
      n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, 
      n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, 
      n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, 
      n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, 
      n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, 
      n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, 
      n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, 
      n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, 
      n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, 
      n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, 
      n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, 
      n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, 
      n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, 
      n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, 
      n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, 
      n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, 
      n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, 
      n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, 
      n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, 
      n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, 
      n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, 
      n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, 
      n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, 
      n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, 
      n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, 
      n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, 
      n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, 
      n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, 
      n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, 
      n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, 
      n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, 
      n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, 
      n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, 
      n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, 
      n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, 
      n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, 
      n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, 
      n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, 
      n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, 
      n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, 
      n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, 
      n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, 
      n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, 
      n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, 
      n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, 
      n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, 
      n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, 
      n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, 
      n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, 
      n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, 
      n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, 
      n17317, n17318, n17319, n17320, n_1000, n_1001, n_1002, n_1003, n_1004, 
      n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, 
      n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT1_reg_31_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => OUT1_31_port
                           , QN => n_1000);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => OUT1_30_port
                           , QN => n_1001);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => OUT1_29_port
                           , QN => n_1002);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => OUT1_28_port
                           , QN => n_1003);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => OUT1_27_port
                           , QN => n_1004);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => OUT1_26_port
                           , QN => n_1005);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => OUT1_25_port
                           , QN => n_1006);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => OUT1_24_port
                           , QN => n_1007);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => OUT1_23_port
                           , QN => n_1008);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => OUT1_22_port
                           , QN => n_1009);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => OUT1_21_port
                           , QN => n_1010);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => OUT1_20_port
                           , QN => n_1011);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => OUT1_19_port
                           , QN => n_1012);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => OUT1_18_port
                           , QN => n_1013);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => OUT1_17_port
                           , QN => n_1014);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => OUT1_16_port
                           , QN => n_1015);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => OUT1_15_port
                           , QN => n_1016);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => OUT1_14_port
                           , QN => n_1017);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => OUT1_13_port
                           , QN => n_1018);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => OUT1_12_port
                           , QN => n_1019);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => OUT1_11_port
                           , QN => n_1020);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => OUT1_10_port
                           , QN => n_1021);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => OUT1_9_port, 
                           QN => n_1022);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => OUT1_8_port, 
                           QN => n_1023);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1024);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1025);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1026);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1027);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1028);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1029);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1030);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1031);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => OUT2_30_port
                           , QN => n_1032);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => OUT2_29_port
                           , QN => n_1033);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => OUT2_28_port
                           , QN => n_1034);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => OUT2_27_port
                           , QN => n_1035);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => OUT2_26_port
                           , QN => n_1036);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => OUT2_25_port
                           , QN => n_1037);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => OUT2_24_port
                           , QN => n_1038);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => OUT2_23_port
                           , QN => n_1039);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => OUT2_22_port
                           , QN => n_1040);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => OUT2_21_port
                           , QN => n_1041);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => OUT2_20_port
                           , QN => n_1042);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => OUT2_19_port
                           , QN => n_1043);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => OUT2_18_port
                           , QN => n_1044);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => OUT2_17_port
                           , QN => n_1045);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => OUT2_16_port
                           , QN => n_1046);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => OUT2_15_port
                           , QN => n_1047);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => OUT2_14_port
                           , QN => n_1048);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => OUT2_13_port
                           , QN => n_1049);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => OUT2_12_port
                           , QN => n_1050);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => OUT2_11_port
                           , QN => n_1051);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => OUT2_10_port
                           , QN => n_1052);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1053);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1054);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1055);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1056);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1057);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1058);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1059);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1060);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1061);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1062);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n_1063, QN => n13690);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n_1064, QN => n13691);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n_1065, QN => n13692);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n_1066, QN => n13693);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n_1067, QN => n13694);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n_1068, QN => n13695);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n_1069, QN => n13696);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n_1070, QN => n13697);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n_1071, QN => n13594);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n_1072, QN => n13595);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n_1073, QN => n13596);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n_1074, QN => n13597);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n_1075, QN => n13598);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n_1076, QN => n13599);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n_1077, QN => n13600);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n_1078, QN => n13601);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n_1079, QN => n13530);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           n_1080, QN => n13531);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n_1081, QN => n13532);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           n_1082, QN => n13533);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n_1083, QN => n13534);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n_1084, QN => n13535);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n_1085, QN => n13536);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n_1086, QN => n13537);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n_1087, QN => n13498);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           n_1088, QN => n13499);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n_1089, QN => n13500);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           n_1090, QN => n13501);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n_1091, QN => n13502);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n_1092, QN => n13503);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n_1093, QN => n13504);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n_1094, QN => n13505);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           n_1095, QN => n13466);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           n_1096, QN => n13467);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           n_1097, QN => n13468);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           n_1098, QN => n13469);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n_1099, QN => n13470);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n_1100, QN => n13471);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n_1101, QN => n13472);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n_1102, QN => n13473);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           n_1103, QN => n13370);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           n_1104, QN => n13371);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           n_1105, QN => n13372);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           n_1106, QN => n13373);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n_1107, QN => n13374);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1108, QN => n13375);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1109, QN => n13376);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1110, QN => n13377);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n_1111, QN => n13338);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n_1112, QN => n13339);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n_1113, QN => n13340);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n_1114, QN => n13341);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n_1115, QN => n13342);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n_1116, QN => n13343);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n_1117, QN => n13344);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n_1118, QN => n13345);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n_1119, QN => n13306);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n_1120, QN => n13307);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n_1121, QN => n13308);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n_1122, QN => n13309);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n_1123, QN => n13310);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n_1124, QN => n13311);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n_1125, QN => n13312);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n_1126, QN => n13313);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n_1127, QN => n13698);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n_1128, QN => n13699);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n_1129, QN => n13700);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n_1130, QN => n13701);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n_1131, QN => n13702);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n_1132, QN => n13703);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n_1133, QN => n13704);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n_1134, QN => n13705);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n_1135, QN => n13706);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n_1136, QN => n13707);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           n_1137, QN => n13708);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           n_1138, QN => n13709);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           n_1139, QN => n13710);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           n_1140, QN => n13711);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           n_1141, QN => n13712);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           n_1142, QN => n13713);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           n_1143, QN => n13714);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           n_1144, QN => n13715);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           n_1145, QN => n13716);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           n_1146, QN => n13717);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           n_1147, QN => n13718);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           n_1148, QN => n13719);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           n_1149, QN => n13720);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           n_1150, QN => n13721);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n_1151, QN => n13602);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n_1152, QN => n13603);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n_1153, QN => n13604);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n_1154, QN => n13605);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n_1155, QN => n13606);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n_1156, QN => n13607);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n_1157, QN => n13608);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n_1158, QN => n13609);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n_1159, QN => n13610);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n_1160, QN => n13611);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           n_1161, QN => n13612);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           n_1162, QN => n13613);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           n_1163, QN => n13614);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           n_1164, QN => n13615);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           n_1165, QN => n13616);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           n_1166, QN => n13617);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           n_1167, QN => n13618);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           n_1168, QN => n13619);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           n_1169, QN => n13620);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           n_1170, QN => n13621);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           n_1171, QN => n13622);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           n_1172, QN => n13623);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           n_1173, QN => n13624);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           n_1174, QN => n13625);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n_1175, QN => n13578);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n_1176, QN => n13579);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n_1177, QN => n13580);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n_1178, QN => n13581);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n_1179, QN => n13582);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n_1180, QN => n13583);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n_1181, QN => n13584);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n_1182, QN => n13585);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n_1183, QN => n13586);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n_1184, QN => n13587);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n_1185, QN => n13588);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n_1186, QN => n13589);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n_1187, QN => n13590);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n_1188, QN => n13591);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n_1189, QN => n13592);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n_1190, QN => n13593);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n_1191, QN => n13538);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n_1192, QN => n13539);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n_1193, QN => n13540);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n_1194, QN => n13541);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n_1195, QN => n13542);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n_1196, QN => n13543);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n_1197, QN => n13544);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n_1198, QN => n13545);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n_1199, QN => n13546);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n_1200, QN => n13547);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n_1201, QN => n13548);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n_1202, QN => n13549);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n_1203, QN => n13550);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n_1204, QN => n13551);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n_1205, QN => n13552);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n_1206, QN => n13553);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n_1207, QN => n13554);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n_1208, QN => n13555);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n_1209, QN => n13556);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           n_1210, QN => n13557);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           n_1211, QN => n13558);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           n_1212, QN => n13559);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           n_1213, QN => n13560);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           n_1214, QN => n13561);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n_1215, QN => n13506);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n_1216, QN => n13507);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n_1217, QN => n13508);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n_1218, QN => n13509);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n_1219, QN => n13510);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n_1220, QN => n13511);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n_1221, QN => n13512);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n_1222, QN => n13513);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n_1223, QN => n13514);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n_1224, QN => n13515);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n_1225, QN => n13516);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n_1226, QN => n13517);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n_1227, QN => n13518);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n_1228, QN => n13519);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n_1229, QN => n13520);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n_1230, QN => n13521);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n_1231, QN => n13522);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n_1232, QN => n13523);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n_1233, QN => n13524);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           n_1234, QN => n13525);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n_1235, QN => n13526);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           n_1236, QN => n13527);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n_1237, QN => n13528);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           n_1238, QN => n13529);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n_1239, QN => n13474);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n_1240, QN => n13475);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n_1241, QN => n13476);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n_1242, QN => n13477);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n_1243, QN => n13478);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n_1244, QN => n13479);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n_1245, QN => n13480);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n_1246, QN => n13481);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n_1247, QN => n13482);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n_1248, QN => n13483);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n_1249, QN => n13484);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n_1250, QN => n13485);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n_1251, QN => n13486);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n_1252, QN => n13487);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n_1253, QN => n13488);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n_1254, QN => n13489);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n_1255, QN => n13490);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n_1256, QN => n13491);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n_1257, QN => n13492);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           n_1258, QN => n13493);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n_1259, QN => n13494);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           n_1260, QN => n13495);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n_1261, QN => n13496);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           n_1262, QN => n13497);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n_1263, QN => n13442);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n_1264, QN => n13443);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n_1265, QN => n13444);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n_1266, QN => n13445);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n_1267, QN => n13446);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n_1268, QN => n13447);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n_1269, QN => n13448);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n_1270, QN => n13449);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n_1271, QN => n13450);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n_1272, QN => n13451);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n_1273, QN => n13452);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n_1274, QN => n13453);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n_1275, QN => n13454);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n_1276, QN => n13455);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n_1277, QN => n13456);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n_1278, QN => n13457);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n_1279, QN => n13458);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n_1280, QN => n13459);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n_1281, QN => n13460);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           n_1282, QN => n13461);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           n_1283, QN => n13462);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           n_1284, QN => n13463);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           n_1285, QN => n13464);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           n_1286, QN => n13465);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n_1287, QN => n13410);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n_1288, QN => n13411);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n_1289, QN => n13412);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n_1290, QN => n13413);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n_1291, QN => n13414);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n_1292, QN => n13415);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n_1293, QN => n13416);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n_1294, QN => n13417);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n_1295, QN => n13418);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n_1296, QN => n13419);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n_1297, QN => n13420);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n_1298, QN => n13421);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n_1299, QN => n13422);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n_1300, QN => n13423);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n_1301, QN => n13424);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n_1302, QN => n13425);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n_1303, QN => n13426);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n_1304, QN => n13427);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           n_1305, QN => n13428);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           n_1306, QN => n13429);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           n_1307, QN => n13430);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           n_1308, QN => n13431);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           n_1309, QN => n13432);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           n_1310, QN => n13433);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1311, QN => n13378);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1312, QN => n13379);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1313, QN => n13380);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1314, QN => n13381);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1315, QN => n13382);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1316, QN => n13383);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1317, QN => n13384);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1318, QN => n13385);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1319, QN => n13386);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1320, QN => n13387);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1321, QN => n13388);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1322, QN => n13389);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1323, QN => n13390);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1324, QN => n13391);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1325, QN => n13392);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1326, QN => n13393);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1327, QN => n13394);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1328, QN => n13395);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1329, QN => n13396);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1330, QN => n13397);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n_1331, QN => n13398);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n_1332, QN => n13399);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n_1333, QN => n13400);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n_1334, QN => n13401);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n_1335, QN => n13346);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n_1336, QN => n13347);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n_1337, QN => n13348);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n_1338, QN => n13349);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n_1339, QN => n13350);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n_1340, QN => n13351);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n_1341, QN => n13352);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n_1342, QN => n13353);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n_1343, QN => n13354);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n_1344, QN => n13355);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n_1345, QN => n13356);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n_1346, QN => n13357);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n_1347, QN => n13358);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n_1348, QN => n13359);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n_1349, QN => n13360);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n_1350, QN => n13361);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n_1351, QN => n13362);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n_1352, QN => n13363);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           n_1353, QN => n13364);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           n_1354, QN => n13365);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           n_1355, QN => n13366);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           n_1356, QN => n13367);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           n_1357, QN => n13368);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           n_1358, QN => n13369);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n_1359, QN => n13314);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n_1360, QN => n13315);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n_1361, QN => n13316);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n_1362, QN => n13317);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n_1363, QN => n13318);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n_1364, QN => n13319);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n_1365, QN => n13320);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n_1366, QN => n13321);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n_1367, QN => n13322);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n_1368, QN => n13323);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n_1369, QN => n13324);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n_1370, QN => n13325);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n_1371, QN => n13326);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n_1372, QN => n13327);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           n_1373, QN => n13328);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           n_1374, QN => n13329);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           n_1375, QN => n13330);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           n_1376, QN => n13331);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           n_1377, QN => n13332);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           n_1378, QN => n13333);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           n_1379, QN => n13334);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           n_1380, QN => n13335);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           n_1381, QN => n13336);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           n_1382, QN => n13337);
   U13672 : NAND3_X1 port map( A1 => n14445, A2 => n14444, A3 => n15143, ZN => 
                           n15135);
   U13673 : NAND3_X1 port map( A1 => n15143, A2 => n14444, A3 => ADD_WR(2), ZN 
                           => n15145);
   U13674 : NAND3_X1 port map( A1 => n15143, A2 => n14445, A3 => ADD_WR(3), ZN 
                           => n15150);
   U13675 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n15143, A3 => ADD_WR(3), 
                           ZN => n15155);
   U13676 : NAND3_X1 port map( A1 => n14445, A2 => n14444, A3 => n15164, ZN => 
                           n15160);
   U13677 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n14444, A3 => n15164, ZN 
                           => n15166);
   U13678 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n14445, A3 => n15164, ZN 
                           => n15171);
   U13679 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n15164, 
                           ZN => n15176);
   U13680 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n16727, A3 => ADD_RD1(1)
                           , ZN => n15220);
   U13684 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n16726, A3 => ADD_RD2(1)
                           , ZN => n15801);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           n_1383, QN => n13722);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           n_1384, QN => n13723);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           n_1385, QN => n13724);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           n_1386, QN => n13725);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           n_1387, QN => n13726);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n_1388, QN => n13727);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n_1389, QN => n13728);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n_1390, QN => n13729);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n_1391, QN => n13730);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n_1392, QN => n13731);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n_1393, QN => n13732);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n_1394, QN => n13733);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n_1395, QN => n13734);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n_1396, QN => n13735);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n_1397, QN => n13736);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n_1398, QN => n13737);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n_1399, QN => n13738);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n_1400, QN => n13739);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           n_1401, QN => n13740);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           n_1402, QN => n13741);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           n_1403, QN => n13742);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           n_1404, QN => n13743);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           n_1405, QN => n13744);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           n_1406, QN => n13745);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           n_1407, QN => n13746);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           n_1408, QN => n13747);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           n_1409, QN => n13748);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           n_1410, QN => n13749);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           n_1411, QN => n13750);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           n_1412, QN => n13751);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           n_1413, QN => n13752);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           n_1414, QN => n13753);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n14845, QN => n13658);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n14846, QN => n13659);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n14847, QN => n13660);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n14848, QN => n13661);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n14849, QN => n13662);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n14850, QN => n13663);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n14851, QN => n13664);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n14852, QN => n13665);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           n14853, QN => n13626);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           n14854, QN => n13627);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           n14855, QN => n13628);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           n14856, QN => n13629);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n14857, QN => n13630);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n14858, QN => n13631);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n14859, QN => n13632);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n14860, QN => n13633);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n14861, QN => n13274);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n14862, QN => n13275);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n14863, QN => n13276);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n14864, QN => n13277);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n14865, QN => n13278);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n14866, QN => n13279);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n14867, QN => n13280);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n14868, QN => n13281);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n14869, QN => n13242);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n14870, QN => n13243);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n14871, QN => n13244);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n14872, QN => n13245);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n14873, QN => n13246);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n14874, QN => n13247);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n14875, QN => n13248);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n14876, QN => n13249);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n14877, QN => n13210);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n14878, QN => n13211);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n14879, QN => n13212);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n14880, QN => n13213);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n14881, QN => n13214);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n14882, QN => n13215);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n14883, QN => n13216);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n14884, QN => n13217);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           n14885, QN => n13082);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           n14886, QN => n13083);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           n14887, QN => n13084);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           n14888, QN => n13085);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           n14889, QN => n13086);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n14890, QN => n13087);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n14891, QN => n13088);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n14892, QN => n13089);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           n14893, QN => n12954);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           n14894, QN => n12955);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           n14895, QN => n12956);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           n14896, QN => n12957);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           n14897, QN => n12958);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           n14898, QN => n12959);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           n14899, QN => n12960);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           n14900, QN => n12961);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => 
                           n14901, QN => n12826);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => 
                           n14902, QN => n12827);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => 
                           n14903, QN => n12828);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => 
                           n14904, QN => n12829);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => 
                           n14905, QN => n12830);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => 
                           n14906, QN => n12831);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => 
                           n14907, QN => n12832);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => 
                           n14908, QN => n12833);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n14909, QN => n13666);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n14910, QN => n13667);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n14911, QN => n13668);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n14912, QN => n13669);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n14913, QN => n13670);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n14914, QN => n13671);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n14915, QN => n13672);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n14916, QN => n13673);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n14917, QN => n13674);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n14918, QN => n13675);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n14919, QN => n13676);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n14920, QN => n13677);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n14921, QN => n13678);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n14922, QN => n13679);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n14923, QN => n13680);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n14924, QN => n13681);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n14925, QN => n13682);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n14926, QN => n13683);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n14927, QN => n13684);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n14928, QN => n13685);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n14929, QN => n13686);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n14930, QN => n13687);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n14931, QN => n13688);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n14932, QN => n13689);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n14933, QN => n13634);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n14934, QN => n13635);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n14935, QN => n13636);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n14936, QN => n13637);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n14937, QN => n13638);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n14938, QN => n13639);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n14939, QN => n13640);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n14940, QN => n13641);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n14941, QN => n13642);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n14942, QN => n13643);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n14943, QN => n13644);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n14944, QN => n13645);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n14945, QN => n13646);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n14946, QN => n13647);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n14947, QN => n13648);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n14948, QN => n13649);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n14949, QN => n13650);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n14950, QN => n13651);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n14951, QN => n13652);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n14952, QN => n13653);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n14953, QN => n13654);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n14954, QN => n13655);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n14955, QN => n13656);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n14956, QN => n13657);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n14957, QN => n13282);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n14958, QN => n13283);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n14959, QN => n13284);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n14960, QN => n13285);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n14961, QN => n13286);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n14962, QN => n13287);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n14963, QN => n13288);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n14964, QN => n13289);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n14965, QN => n13290);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n14966, QN => n13291);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n14967, QN => n13292);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n14968, QN => n13293);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n14969, QN => n13294);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n14970, QN => n13295);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n14971, QN => n13296);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n14972, QN => n13297);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n14973, QN => n13298);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n14974, QN => n13299);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n14975, QN => n13300);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           n14976, QN => n13301);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           n14977, QN => n13302);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           n14978, QN => n13303);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           n14979, QN => n13304);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           n14980, QN => n13305);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n14981, QN => n13250);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n14982, QN => n13251);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n14983, QN => n13252);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n14984, QN => n13253);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n14985, QN => n13254);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n14986, QN => n13255);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n14987, QN => n13256);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n14988, QN => n13257);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n14989, QN => n13258);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n14990, QN => n13259);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n14991, QN => n13260);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n14992, QN => n13261);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n14993, QN => n13262);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n14994, QN => n13263);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           n14995, QN => n13264);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           n14996, QN => n13265);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           n14997, QN => n13266);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           n14998, QN => n13267);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           n14999, QN => n13268);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           n15000, QN => n13269);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           n15001, QN => n13270);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           n15002, QN => n13271);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           n15003, QN => n13272);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           n15004, QN => n13273);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n15005, QN => n13218);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n15006, QN => n13219);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n15007, QN => n13220);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n15008, QN => n13221);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n15009, QN => n13222);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n15010, QN => n13223);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n15011, QN => n13224);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n15012, QN => n13225);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n15013, QN => n13226);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n15014, QN => n13227);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n15015, QN => n13228);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n15016, QN => n13229);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n15017, QN => n13230);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n15018, QN => n13231);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n15019, QN => n13232);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n15020, QN => n13233);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n15021, QN => n13234);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n15022, QN => n13235);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n15023, QN => n13236);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n15024, QN => n13237);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n15025, QN => n13238);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n15026, QN => n13239);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n15027, QN => n13240);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n15028, QN => n13241);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n15029, QN => n13090);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n15030, QN => n13091);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n15031, QN => n13092);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n15032, QN => n13093);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n15033, QN => n13094);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n15034, QN => n13095);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n15035, QN => n13096);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n15036, QN => n13097);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n15037, QN => n13098);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n15038, QN => n13099);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n15039, QN => n13100);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n15040, QN => n13101);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n15041, QN => n13102);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n15042, QN => n13103);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n15043, QN => n13104);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n15044, QN => n13105);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n15045, QN => n13106);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n15046, QN => n13107);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           n15047, QN => n13108);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           n15048, QN => n13109);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           n15049, QN => n13110);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           n15050, QN => n13111);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           n15051, QN => n13112);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           n15052, QN => n13113);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           n15053, QN => n12962);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           n15054, QN => n12963);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           n15055, QN => n12964);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           n15056, QN => n12965);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           n15057, QN => n12966);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           n15058, QN => n12967);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           n15059, QN => n12968);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           n15060, QN => n12969);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           n15061, QN => n12970);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           n15062, QN => n12971);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           n15063, QN => n12972);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           n15064, QN => n12973);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           n15065, QN => n12974);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           n15066, QN => n12975);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => n15067
                           , QN => n12976);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => n15068
                           , QN => n12977);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => n15069
                           , QN => n12978);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => n15070
                           , QN => n12979);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => n15071
                           , QN => n12980);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n15072
                           , QN => n12981);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => n15073
                           , QN => n12982);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => n15074
                           , QN => n12983);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => n15075
                           , QN => n12984);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => n15076
                           , QN => n12985);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => 
                           n15077, QN => n12834);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => 
                           n15078, QN => n12835);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => 
                           n15079, QN => n12836);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => 
                           n15080, QN => n12837);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => 
                           n15081, QN => n12838);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => 
                           n15082, QN => n12839);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => 
                           n15083, QN => n12840);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => 
                           n15084, QN => n12841);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => 
                           n15085, QN => n12842);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => 
                           n15086, QN => n12843);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => 
                           n15087, QN => n12844);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => 
                           n15088, QN => n12845);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => 
                           n15089, QN => n12846);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => 
                           n15090, QN => n12847);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => n15091
                           , QN => n12848);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => n15092
                           , QN => n12849);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => n15093
                           , QN => n12850);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => n15094
                           , QN => n12851);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => n15095
                           , QN => n12852);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => n15096
                           , QN => n12853);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => n15097
                           , QN => n12854);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => n15098
                           , QN => n12855);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => n15099
                           , QN => n12856);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => n15100
                           , QN => n12857);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           n_1415, QN => n13562);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           n_1416, QN => n13563);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           n_1417, QN => n13564);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           n_1418, QN => n13565);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n_1419, QN => n13566);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n_1420, QN => n13567);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n_1421, QN => n13568);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n_1422, QN => n13569);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1423, QN => n13402);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1424, QN => n13403);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1425, QN => n13404);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1426, QN => n13405);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n_1427, QN => n13406);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n_1428, QN => n13407);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n_1429, QN => n13408);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n_1430, QN => n13409);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           n_1431, QN => n13434);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           n_1432, QN => n13435);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           n_1433, QN => n13436);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           n_1434, QN => n13437);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n_1435, QN => n13438);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n_1436, QN => n13439);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n_1437, QN => n13440);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n_1438, QN => n13441);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n_1439, QN => n13570);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n_1440, QN => n13571);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n_1441, QN => n13572);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n_1442, QN => n13573);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n_1443, QN => n13574);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n_1444, QN => n13575);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n_1445, QN => n13576);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n_1446, QN => n13577);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           n_1447, QN => n15101);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           n_1448, QN => n14814);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           n_1449, QN => n14815);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           n_1450, QN => n14816);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n_1451, QN => n14817);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n_1452, QN => n14818);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n_1453, QN => n14819);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n_1454, QN => n14820);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => 
                           n_1455, QN => n14622);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => 
                           n_1456, QN => n14623);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => 
                           n_1457, QN => n14624);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => 
                           n_1458, QN => n14625);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => 
                           n_1459, QN => n14626);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           n_1460, QN => n14627);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           n_1461, QN => n14628);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           n_1462, QN => n14629);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           n_1463, QN => n14782);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           n_1464, QN => n14783);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n_1465, QN => n14784);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n_1466, QN => n14785);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n_1467, QN => n14786);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n_1468, QN => n14787);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n_1469, QN => n14788);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           n_1470, QN => n14789);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => 
                           n_1471, QN => n14590);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => 
                           n_1472, QN => n14591);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => 
                           n_1473, QN => n14592);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => 
                           n_1474, QN => n14593);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => 
                           n_1475, QN => n14594);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => 
                           n_1476, QN => n14595);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => 
                           n_1477, QN => n14596);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => 
                           n_1478, QN => n14597);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           n_1479, QN => n14750);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           n_1480, QN => n14751);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           n_1481, QN => n14752);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           n_1482, QN => n14753);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n_1483, QN => n14754);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n_1484, QN => n14755);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n_1485, QN => n14756);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n_1486, QN => n14757);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => 
                           n_1487, QN => n14558);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => 
                           n_1488, QN => n14559);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => 
                           n_1489, QN => n14560);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => 
                           n_1490, QN => n14561);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => 
                           n_1491, QN => n14562);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => 
                           n_1492, QN => n14563);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => 
                           n_1493, QN => n14564);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => 
                           n_1494, QN => n14565);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n_1495, QN => n14821);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n_1496, QN => n14822);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n_1497, QN => n14823);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n_1498, QN => n14824);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n_1499, QN => n14825);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n_1500, QN => n14826);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n_1501, QN => n14827);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n_1502, QN => n14828);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n_1503, QN => n14829);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n_1504, QN => n14830);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n_1505, QN => n14831);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n_1506, QN => n14832);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n_1507, QN => n14833);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n_1508, QN => n14834);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n_1509, QN => n14835);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n_1510, QN => n14836);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n_1511, QN => n14837);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n_1512, QN => n14838);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           n_1513, QN => n14839);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           n_1514, QN => n14840);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           n_1515, QN => n14841);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           n_1516, QN => n14842);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           n_1517, QN => n14843);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           n_1518, QN => n14844);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           n_1519, QN => n14630);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           n_1520, QN => n14631);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           n_1521, QN => n14632);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           n_1522, QN => n14633);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           n_1523, QN => n14634);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           n_1524, QN => n14635);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           n_1525, QN => n14636);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           n_1526, QN => n14637);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           n_1527, QN => n14638);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           n_1528, QN => n14639);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           n_1529, QN => n14640);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           n_1530, QN => n14641);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           n_1531, QN => n14642);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           n_1532, QN => n14643);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => n_1533
                           , QN => n14644);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => n_1534
                           , QN => n14645);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => n_1535
                           , QN => n14646);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => n_1536
                           , QN => n14647);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => n_1537
                           , QN => n14648);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n_1538
                           , QN => n14649);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => n_1539
                           , QN => n14650);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => n_1540
                           , QN => n14651);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => n_1541
                           , QN => n14652);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => n_1542
                           , QN => n14653);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           n_1543, QN => n14790);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           n_1544, QN => n14791);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           n_1545, QN => n14792);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           n_1546, QN => n14793);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           n_1547, QN => n14794);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           n_1548, QN => n14795);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           n_1549, QN => n14796);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           n_1550, QN => n14797);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           n_1551, QN => n14798);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n_1552, QN => n14799);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           n_1553, QN => n14800);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           n_1554, QN => n14801);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           n_1555, QN => n14802);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           n_1556, QN => n14803);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           n_1557, QN => n14804);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           n_1558, QN => n14805);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           n_1559, QN => n14806);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           n_1560, QN => n14807);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           n_1561, QN => n14808);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           n_1562, QN => n14809);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           n_1563, QN => n14810);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           n_1564, QN => n14811);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           n_1565, QN => n14812);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           n_1566, QN => n14813);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => 
                           n_1567, QN => n14598);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => 
                           n_1568, QN => n14599);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => 
                           n_1569, QN => n14600);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => 
                           n_1570, QN => n14601);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => 
                           n_1571, QN => n14602);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => 
                           n_1572, QN => n14603);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => 
                           n_1573, QN => n14604);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => 
                           n_1574, QN => n14605);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => 
                           n_1575, QN => n14606);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => 
                           n_1576, QN => n14607);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => 
                           n_1577, QN => n14608);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => 
                           n_1578, QN => n14609);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => 
                           n_1579, QN => n14610);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => 
                           n_1580, QN => n14611);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => n_1581
                           , QN => n14612);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => n_1582
                           , QN => n14613);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => n_1583
                           , QN => n14614);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => n_1584
                           , QN => n14615);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => n_1585
                           , QN => n14616);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n_1586
                           , QN => n14617);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => n_1587
                           , QN => n14618);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => n_1588
                           , QN => n14619);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => n_1589
                           , QN => n14620);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => n_1590
                           , QN => n14621);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           n_1591, QN => n14686);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           n_1592, QN => n14687);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           n_1593, QN => n14688);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           n_1594, QN => n14689);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           n_1595, QN => n14690);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n_1596, QN => n14691);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n_1597, QN => n14692);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           n_1598, QN => n14693);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n_1599, QN => n14758);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n_1600, QN => n14759);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n_1601, QN => n14760);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n_1602, QN => n14761);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n_1603, QN => n14762);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n_1604, QN => n14763);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n_1605, QN => n14764);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n_1606, QN => n14765);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n_1607, QN => n14766);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n_1608, QN => n14767);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           n_1609, QN => n14768);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           n_1610, QN => n14769);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           n_1611, QN => n14770);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           n_1612, QN => n14771);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           n_1613, QN => n14772);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           n_1614, QN => n14773);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           n_1615, QN => n14774);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           n_1616, QN => n14775);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           n_1617, QN => n14776);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           n_1618, QN => n14777);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           n_1619, QN => n14778);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           n_1620, QN => n14779);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           n_1621, QN => n14780);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           n_1622, QN => n14781);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => 
                           n_1623, QN => n14566);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => 
                           n_1624, QN => n14567);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => 
                           n_1625, QN => n14568);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => 
                           n_1626, QN => n14569);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => 
                           n_1627, QN => n14570);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => 
                           n_1628, QN => n14571);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => 
                           n_1629, QN => n14572);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => 
                           n_1630, QN => n14573);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => 
                           n_1631, QN => n14574);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => 
                           n_1632, QN => n14575);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => 
                           n_1633, QN => n14576);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => 
                           n_1634, QN => n14577);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => 
                           n_1635, QN => n14578);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => 
                           n_1636, QN => n14579);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => n_1637
                           , QN => n14580);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => n_1638
                           , QN => n14581);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => n_1639
                           , QN => n14582);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => n_1640
                           , QN => n14583);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => n_1641
                           , QN => n14584);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => n_1642
                           , QN => n14585);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => n_1643
                           , QN => n14586);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => n_1644
                           , QN => n14587);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => n_1645
                           , QN => n14588);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => n_1646
                           , QN => n14589);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           n_1647, QN => n14694);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           n_1648, QN => n14695);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           n_1649, QN => n14696);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           n_1650, QN => n14697);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           n_1651, QN => n14698);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           n_1652, QN => n14699);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           n_1653, QN => n14700);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           n_1654, QN => n14701);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           n_1655, QN => n14702);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           n_1656, QN => n14703);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           n_1657, QN => n14704);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           n_1658, QN => n14705);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           n_1659, QN => n14706);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           n_1660, QN => n14707);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => n_1661
                           , QN => n14708);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => n_1662
                           , QN => n14709);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => n_1663
                           , QN => n14710);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => n_1664
                           , QN => n14711);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => n_1665
                           , QN => n14712);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n_1666
                           , QN => n14713);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => n_1667
                           , QN => n14714);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => n_1668
                           , QN => n14715);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => n_1669
                           , QN => n14716);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => n_1670
                           , QN => n14717);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2331, CK => CLK, Q => 
                           n16429, QN => n14494);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2330, CK => CLK, Q => 
                           n16428, QN => n14495);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2329, CK => CLK, Q => 
                           n16427, QN => n14496);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2328, CK => CLK, Q => 
                           n16426, QN => n14497);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2327, CK => CLK, Q => 
                           n16425, QN => n14498);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2326, CK => CLK, Q => 
                           n16424, QN => n14499);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2325, CK => CLK, Q => 
                           n16423, QN => n14500);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2324, CK => CLK, Q => 
                           n16422, QN => n14501);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2323, CK => CLK, Q => 
                           n16557, QN => n14502);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2322, CK => CLK, Q => 
                           n16556, QN => n14503);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2321, CK => CLK, Q => 
                           n16555, QN => n14504);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2320, CK => CLK, Q => 
                           n16554, QN => n14505);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2319, CK => CLK, Q => 
                           n16553, QN => n14506);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2318, CK => CLK, Q => 
                           n16552, QN => n14507);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2317, CK => CLK, Q => 
                           n16551, QN => n14508);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2316, CK => CLK, Q => 
                           n16550, QN => n14509);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2315, CK => CLK, Q => 
                           n16549, QN => n14510);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2314, CK => CLK, Q => 
                           n16548, QN => n14511);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2313, CK => CLK, Q => 
                           n16547, QN => n14512);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2312, CK => CLK, Q => 
                           n16546, QN => n14513);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2311, CK => CLK, Q => 
                           n16545, QN => n14514);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2310, CK => CLK, Q => 
                           n16544, QN => n14515);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2309, CK => CLK, Q => n16543
                           , QN => n14516);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2308, CK => CLK, Q => n16542
                           , QN => n14517);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2307, CK => CLK, Q => n16541
                           , QN => n14518);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2306, CK => CLK, Q => n16540
                           , QN => n14519);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2305, CK => CLK, Q => n16539
                           , QN => n14520);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2304, CK => CLK, Q => n16538
                           , QN => n14521);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2303, CK => CLK, Q => n16537
                           , QN => n14522);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2302, CK => CLK, Q => n16536
                           , QN => n14523);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2301, CK => CLK, Q => n16535
                           , QN => n14524);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2300, CK => CLK, Q => n16534
                           , QN => n14525);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           n16373, QN => n14718);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           n16372, QN => n14719);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           n16371, QN => n14720);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           n16370, QN => n14721);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           n16369, QN => n14722);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           n16368, QN => n14723);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           n16367, QN => n14724);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           n16366, QN => n14725);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           n16677, QN => n14726);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           n16676, QN => n14727);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           n16675, QN => n14728);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           n16674, QN => n14729);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           n16673, QN => n14730);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           n16672, QN => n14731);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           n16671, QN => n14732);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           n16670, QN => n14733);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           n16669, QN => n14734);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           n16668, QN => n14735);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           n16667, QN => n14736);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           n16666, QN => n14737);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           n16665, QN => n14738);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           n16664, QN => n14739);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           n16663, QN => n14740);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           n16662, QN => n14741);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           n16661, QN => n14742);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           n16660, QN => n14743);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           n16659, QN => n14744);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           n16658, QN => n14745);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           n16657, QN => n14746);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           n16656, QN => n14747);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           n16655, QN => n14748);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           n16654, QN => n14749);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           n16389, QN => n14654);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           n16388, QN => n14655);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           n16387, QN => n14656);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           n16386, QN => n14657);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           n16385, QN => n14658);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           n16384, QN => n14659);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           n16383, QN => n14660);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           n16382, QN => n14661);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2363, CK => CLK, Q => 
                           n16437, QN => n14462);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2362, CK => CLK, Q => 
                           n16436, QN => n14463);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2361, CK => CLK, Q => 
                           n16435, QN => n14464);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2360, CK => CLK, Q => 
                           n16434, QN => n14465);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2359, CK => CLK, Q => 
                           n16433, QN => n14466);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2358, CK => CLK, Q => 
                           n16432, QN => n14467);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2357, CK => CLK, Q => 
                           n16431, QN => n14468);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2356, CK => CLK, Q => 
                           n16430, QN => n14469);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2299, CK => CLK, Q => 
                           n16421, QN => n14526);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2298, CK => CLK, Q => 
                           n16420, QN => n14527);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2297, CK => CLK, Q => 
                           n16419, QN => n14528);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2296, CK => CLK, Q => 
                           n16418, QN => n14529);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => 
                           n16417, QN => n14530);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => 
                           n16416, QN => n14531);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => 
                           n16415, QN => n14532);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => 
                           n16414, QN => n14533);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           n16725, QN => n14662);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           n16724, QN => n14663);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           n16723, QN => n14664);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           n16722, QN => n14665);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           n16721, QN => n14666);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           n16720, QN => n14667);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           n16719, QN => n14668);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           n16718, QN => n14669);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           n16717, QN => n14670);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           n16716, QN => n14671);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           n16715, QN => n14672);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           n16714, QN => n14673);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           n16713, QN => n14674);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           n16712, QN => n14675);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => n16711
                           , QN => n14676);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => n16710
                           , QN => n14677);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => n16709
                           , QN => n14678);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => n16708
                           , QN => n14679);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => n16707
                           , QN => n14680);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n16706
                           , QN => n14681);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n16705
                           , QN => n14682);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n16704
                           , QN => n14683);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => n16703
                           , QN => n14684);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => n16702
                           , QN => n14685);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2355, CK => CLK, Q => 
                           n16581, QN => n14470);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2354, CK => CLK, Q => 
                           n16580, QN => n14471);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2353, CK => CLK, Q => 
                           n16579, QN => n14472);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2352, CK => CLK, Q => 
                           n16578, QN => n14473);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2351, CK => CLK, Q => 
                           n16577, QN => n14474);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2350, CK => CLK, Q => 
                           n16576, QN => n14475);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2349, CK => CLK, Q => 
                           n16575, QN => n14476);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2348, CK => CLK, Q => 
                           n16574, QN => n14477);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2347, CK => CLK, Q => 
                           n16573, QN => n14478);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2346, CK => CLK, Q => 
                           n16572, QN => n14479);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2345, CK => CLK, Q => 
                           n16571, QN => n14480);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2344, CK => CLK, Q => 
                           n16570, QN => n14481);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2343, CK => CLK, Q => 
                           n16569, QN => n14482);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2342, CK => CLK, Q => 
                           n16568, QN => n14483);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2341, CK => CLK, Q => n16567
                           , QN => n14484);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2340, CK => CLK, Q => n16566
                           , QN => n14485);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2339, CK => CLK, Q => n16565
                           , QN => n14486);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2338, CK => CLK, Q => n16564
                           , QN => n14487);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2337, CK => CLK, Q => n16563
                           , QN => n14488);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2336, CK => CLK, Q => n16562
                           , QN => n14489);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2335, CK => CLK, Q => n16561
                           , QN => n14490);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2334, CK => CLK, Q => n16560
                           , QN => n14491);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2333, CK => CLK, Q => n16559
                           , QN => n14492);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2332, CK => CLK, Q => n16558
                           , QN => n14493);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => 
                           n16533, QN => n14534);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => 
                           n16532, QN => n14535);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => 
                           n16531, QN => n14536);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => 
                           n16530, QN => n14537);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => 
                           n16529, QN => n14538);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => 
                           n16528, QN => n14539);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => 
                           n16527, QN => n14540);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => 
                           n16526, QN => n14541);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => 
                           n16525, QN => n14542);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => 
                           n16524, QN => n14543);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => 
                           n16523, QN => n14544);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => 
                           n16522, QN => n14545);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => 
                           n16521, QN => n14546);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => 
                           n16520, QN => n14547);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => n16519
                           , QN => n14548);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => n16518
                           , QN => n14549);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => n16517
                           , QN => n14550);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => n16516
                           , QN => n14551);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => n16515
                           , QN => n14552);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => n16514
                           , QN => n14553);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => n16513
                           , QN => n14554);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => n16512
                           , QN => n14555);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => n16511
                           , QN => n14556);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => n16510
                           , QN => n14557);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => OUT2_31_port
                           , QN => n_1671);
   U13688 : NOR3_X1 port map( A1 => n16754, A2 => ADD_RD2(0), A3 => n14461, ZN 
                           => n16331);
   U13689 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n16754,
                           ZN => n16330);
   U13690 : NOR3_X1 port map( A1 => n16847, A2 => ADD_RD1(0), A3 => n14454, ZN 
                           => n15750);
   U13691 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n16847,
                           ZN => n15749);
   U13692 : INV_X1 port map( A => n17061, ZN => n17054);
   U13693 : INV_X1 port map( A => n17298, ZN => n17291);
   U13694 : INV_X1 port map( A => n17178, ZN => n17171);
   U13695 : INV_X1 port map( A => n17142, ZN => n17135);
   U13696 : INV_X1 port map( A => n17106, ZN => n17099);
   U13697 : INV_X1 port map( A => n17070, ZN => n17063);
   U13698 : INV_X1 port map( A => n17052, ZN => n17045);
   U13699 : INV_X1 port map( A => n17043, ZN => n17036);
   U13700 : INV_X1 port map( A => n17034, ZN => n17027);
   U13701 : INV_X1 port map( A => n17025, ZN => n17018);
   U13702 : INV_X1 port map( A => n17016, ZN => n17009);
   U13703 : INV_X1 port map( A => n17007, ZN => n17000);
   U13704 : INV_X1 port map( A => n16998, ZN => n16991);
   U13705 : INV_X1 port map( A => n16989, ZN => n16982);
   U13706 : INV_X1 port map( A => n16980, ZN => n16973);
   U13707 : INV_X1 port map( A => n16971, ZN => n16964);
   U13708 : INV_X1 port map( A => n16962, ZN => n16955);
   U13709 : INV_X1 port map( A => n16953, ZN => n16946);
   U13710 : INV_X1 port map( A => n16944, ZN => n16937);
   U13711 : INV_X1 port map( A => n16935, ZN => n16928);
   U13712 : INV_X1 port map( A => n17079, ZN => n17072);
   U13713 : INV_X1 port map( A => n17088, ZN => n17081);
   U13714 : INV_X1 port map( A => n17097, ZN => n17090);
   U13715 : INV_X1 port map( A => n17115, ZN => n17108);
   U13716 : INV_X1 port map( A => n17124, ZN => n17117);
   U13717 : INV_X1 port map( A => n17133, ZN => n17126);
   U13718 : INV_X1 port map( A => n17151, ZN => n17144);
   U13719 : INV_X1 port map( A => n17160, ZN => n17153);
   U13720 : INV_X1 port map( A => n17169, ZN => n17162);
   U13721 : INV_X1 port map( A => n17187, ZN => n17180);
   U13722 : INV_X1 port map( A => n17196, ZN => n17189);
   U13723 : BUF_X1 port map( A => n17062, Z => n17055);
   U13724 : BUF_X1 port map( A => n17062, Z => n17056);
   U13725 : BUF_X1 port map( A => n17062, Z => n17057);
   U13726 : BUF_X1 port map( A => n17062, Z => n17058);
   U13727 : BUF_X1 port map( A => n17062, Z => n17059);
   U13728 : BUF_X1 port map( A => n17062, Z => n17060);
   U13729 : BUF_X1 port map( A => n17299, Z => n17292);
   U13730 : BUF_X1 port map( A => n17299, Z => n17293);
   U13731 : BUF_X1 port map( A => n17299, Z => n17294);
   U13732 : BUF_X1 port map( A => n17299, Z => n17295);
   U13733 : BUF_X1 port map( A => n17299, Z => n17296);
   U13734 : BUF_X1 port map( A => n17299, Z => n17297);
   U13735 : BUF_X1 port map( A => n17062, Z => n17061);
   U13736 : BUF_X1 port map( A => n17299, Z => n17298);
   U13737 : BUF_X1 port map( A => n16927, Z => n16919);
   U13738 : BUF_X1 port map( A => n16927, Z => n16920);
   U13739 : BUF_X1 port map( A => n16927, Z => n16921);
   U13740 : BUF_X1 port map( A => n16927, Z => n16922);
   U13741 : BUF_X1 port map( A => n16927, Z => n16923);
   U13742 : BUF_X1 port map( A => n16927, Z => n16924);
   U13743 : BUF_X1 port map( A => n16924, Z => n16925);
   U13744 : BUF_X1 port map( A => n16919, Z => n16926);
   U13745 : BUF_X1 port map( A => n15786, Z => n16780);
   U13746 : BUF_X1 port map( A => n15786, Z => n16781);
   U13747 : BUF_X1 port map( A => n15205, Z => n16873);
   U13748 : BUF_X1 port map( A => n15205, Z => n16874);
   U13749 : BUF_X1 port map( A => n14457, Z => n17306);
   U13750 : BUF_X1 port map( A => n14457, Z => n17307);
   U13751 : BUF_X1 port map( A => n14450, Z => n17312);
   U13752 : BUF_X1 port map( A => n14450, Z => n17313);
   U13753 : BUF_X1 port map( A => n15787, Z => n16777);
   U13754 : BUF_X1 port map( A => n15787, Z => n16778);
   U13755 : BUF_X1 port map( A => n15206, Z => n16870);
   U13756 : BUF_X1 port map( A => n15206, Z => n16871);
   U13757 : BUF_X1 port map( A => n14458, Z => n17303);
   U13758 : BUF_X1 port map( A => n14458, Z => n17304);
   U13759 : BUF_X1 port map( A => n14451, Z => n17309);
   U13760 : BUF_X1 port map( A => n14451, Z => n17310);
   U13761 : BUF_X1 port map( A => n15789, Z => n16771);
   U13762 : BUF_X1 port map( A => n15789, Z => n16772);
   U13763 : BUF_X1 port map( A => n15208, Z => n16864);
   U13764 : BUF_X1 port map( A => n15208, Z => n16865);
   U13765 : BUF_X1 port map( A => n15779, Z => n16792);
   U13766 : BUF_X1 port map( A => n15779, Z => n16793);
   U13767 : BUF_X1 port map( A => n15198, Z => n16885);
   U13768 : BUF_X1 port map( A => n15198, Z => n16886);
   U13769 : BUF_X1 port map( A => n15783, Z => n16783);
   U13770 : BUF_X1 port map( A => n15783, Z => n16784);
   U13771 : BUF_X1 port map( A => n15202, Z => n16876);
   U13772 : BUF_X1 port map( A => n15202, Z => n16877);
   U13773 : BUF_X1 port map( A => n15793, Z => n16762);
   U13774 : BUF_X1 port map( A => n15793, Z => n16763);
   U13775 : BUF_X1 port map( A => n15212, Z => n16855);
   U13776 : BUF_X1 port map( A => n15212, Z => n16856);
   U13777 : BUF_X1 port map( A => n15791, Z => n16768);
   U13778 : BUF_X1 port map( A => n15781, Z => n16789);
   U13779 : BUF_X1 port map( A => n15791, Z => n16769);
   U13780 : BUF_X1 port map( A => n15781, Z => n16790);
   U13781 : BUF_X1 port map( A => n15210, Z => n16861);
   U13782 : BUF_X1 port map( A => n15200, Z => n16882);
   U13783 : BUF_X1 port map( A => n15210, Z => n16862);
   U13784 : BUF_X1 port map( A => n15200, Z => n16883);
   U13785 : BUF_X1 port map( A => n15797, Z => n16751);
   U13786 : BUF_X1 port map( A => n15797, Z => n16752);
   U13787 : BUF_X1 port map( A => n15216, Z => n16844);
   U13788 : BUF_X1 port map( A => n15216, Z => n16845);
   U13789 : BUF_X1 port map( A => n15788, Z => n16774);
   U13790 : BUF_X1 port map( A => n15788, Z => n16775);
   U13791 : BUF_X1 port map( A => n15207, Z => n16867);
   U13792 : BUF_X1 port map( A => n15207, Z => n16868);
   U13793 : BUF_X1 port map( A => n15778, Z => n16795);
   U13794 : BUF_X1 port map( A => n15778, Z => n16796);
   U13795 : BUF_X1 port map( A => n15197, Z => n16888);
   U13796 : BUF_X1 port map( A => n15197, Z => n16889);
   U13797 : BUF_X1 port map( A => n15771, Z => n16816);
   U13798 : BUF_X1 port map( A => n15774, Z => n16807);
   U13799 : BUF_X1 port map( A => n15777, Z => n16798);
   U13800 : BUF_X1 port map( A => n15771, Z => n16817);
   U13801 : BUF_X1 port map( A => n15774, Z => n16808);
   U13802 : BUF_X1 port map( A => n15777, Z => n16799);
   U13803 : BUF_X1 port map( A => n15190, Z => n16909);
   U13804 : BUF_X1 port map( A => n15193, Z => n16900);
   U13805 : BUF_X1 port map( A => n15196, Z => n16891);
   U13806 : BUF_X1 port map( A => n15190, Z => n16910);
   U13807 : BUF_X1 port map( A => n15193, Z => n16901);
   U13808 : BUF_X1 port map( A => n15196, Z => n16892);
   U13809 : BUF_X1 port map( A => n15786, Z => n16782);
   U13810 : BUF_X1 port map( A => n15205, Z => n16875);
   U13811 : BUF_X1 port map( A => n14457, Z => n17308);
   U13812 : BUF_X1 port map( A => n14450, Z => n17314);
   U13813 : BUF_X1 port map( A => n15794, Z => n16760);
   U13814 : BUF_X1 port map( A => n15794, Z => n16759);
   U13815 : BUF_X1 port map( A => n15213, Z => n16853);
   U13816 : BUF_X1 port map( A => n15213, Z => n16852);
   U13817 : BUF_X1 port map( A => n15769, Z => n16822);
   U13818 : BUF_X1 port map( A => n15772, Z => n16813);
   U13819 : BUF_X1 port map( A => n15775, Z => n16804);
   U13820 : BUF_X1 port map( A => n15769, Z => n16823);
   U13821 : BUF_X1 port map( A => n15772, Z => n16814);
   U13822 : BUF_X1 port map( A => n15775, Z => n16805);
   U13823 : BUF_X1 port map( A => n15188, Z => n16915);
   U13824 : BUF_X1 port map( A => n15191, Z => n16906);
   U13825 : BUF_X1 port map( A => n15194, Z => n16897);
   U13826 : BUF_X1 port map( A => n15188, Z => n16916);
   U13827 : BUF_X1 port map( A => n15191, Z => n16907);
   U13828 : BUF_X1 port map( A => n15194, Z => n16898);
   U13829 : BUF_X1 port map( A => n15770, Z => n16819);
   U13830 : BUF_X1 port map( A => n15773, Z => n16810);
   U13831 : BUF_X1 port map( A => n15776, Z => n16801);
   U13832 : BUF_X1 port map( A => n15770, Z => n16820);
   U13833 : BUF_X1 port map( A => n15773, Z => n16811);
   U13834 : BUF_X1 port map( A => n15776, Z => n16802);
   U13835 : BUF_X1 port map( A => n15189, Z => n16912);
   U13836 : BUF_X1 port map( A => n15192, Z => n16903);
   U13837 : BUF_X1 port map( A => n15195, Z => n16894);
   U13838 : BUF_X1 port map( A => n15189, Z => n16913);
   U13839 : BUF_X1 port map( A => n15192, Z => n16904);
   U13840 : BUF_X1 port map( A => n15195, Z => n16895);
   U13841 : BUF_X1 port map( A => n15787, Z => n16779);
   U13842 : BUF_X1 port map( A => n15206, Z => n16872);
   U13843 : BUF_X1 port map( A => n14458, Z => n17305);
   U13844 : BUF_X1 port map( A => n14451, Z => n17311);
   U13845 : BUF_X1 port map( A => n15792, Z => n16766);
   U13846 : BUF_X1 port map( A => n15782, Z => n16787);
   U13847 : BUF_X1 port map( A => n15792, Z => n16765);
   U13848 : BUF_X1 port map( A => n15782, Z => n16786);
   U13849 : BUF_X1 port map( A => n15211, Z => n16859);
   U13850 : BUF_X1 port map( A => n15201, Z => n16880);
   U13851 : BUF_X1 port map( A => n15211, Z => n16858);
   U13852 : BUF_X1 port map( A => n15201, Z => n16879);
   U13853 : BUF_X1 port map( A => n15795, Z => n16757);
   U13854 : BUF_X1 port map( A => n15795, Z => n16756);
   U13855 : BUF_X1 port map( A => n15214, Z => n16850);
   U13856 : BUF_X1 port map( A => n15214, Z => n16849);
   U13857 : BUF_X1 port map( A => n15789, Z => n16773);
   U13858 : BUF_X1 port map( A => n15208, Z => n16866);
   U13859 : BUF_X1 port map( A => n15779, Z => n16794);
   U13860 : BUF_X1 port map( A => n15198, Z => n16887);
   U13861 : BUF_X1 port map( A => n15783, Z => n16785);
   U13862 : BUF_X1 port map( A => n15202, Z => n16878);
   U13863 : BUF_X1 port map( A => n15793, Z => n16764);
   U13864 : BUF_X1 port map( A => n15212, Z => n16857);
   U13865 : BUF_X1 port map( A => n15791, Z => n16770);
   U13866 : BUF_X1 port map( A => n15781, Z => n16791);
   U13867 : BUF_X1 port map( A => n15210, Z => n16863);
   U13868 : BUF_X1 port map( A => n15200, Z => n16884);
   U13869 : BUF_X1 port map( A => n15797, Z => n16753);
   U13870 : BUF_X1 port map( A => n15216, Z => n16846);
   U13871 : BUF_X1 port map( A => n15788, Z => n16776);
   U13872 : BUF_X1 port map( A => n15207, Z => n16869);
   U13873 : BUF_X1 port map( A => n15778, Z => n16797);
   U13874 : BUF_X1 port map( A => n15197, Z => n16890);
   U13875 : BUF_X1 port map( A => n15771, Z => n16818);
   U13876 : BUF_X1 port map( A => n15774, Z => n16809);
   U13877 : BUF_X1 port map( A => n15777, Z => n16800);
   U13878 : BUF_X1 port map( A => n15190, Z => n16911);
   U13879 : BUF_X1 port map( A => n15193, Z => n16902);
   U13880 : BUF_X1 port map( A => n15196, Z => n16893);
   U13881 : BUF_X1 port map( A => n15794, Z => n16761);
   U13882 : BUF_X1 port map( A => n15213, Z => n16854);
   U13883 : BUF_X1 port map( A => n15769, Z => n16824);
   U13884 : BUF_X1 port map( A => n15772, Z => n16815);
   U13885 : BUF_X1 port map( A => n15775, Z => n16806);
   U13886 : BUF_X1 port map( A => n15188, Z => n16917);
   U13887 : BUF_X1 port map( A => n15191, Z => n16908);
   U13888 : BUF_X1 port map( A => n15194, Z => n16899);
   U13889 : BUF_X1 port map( A => n15770, Z => n16821);
   U13890 : BUF_X1 port map( A => n15773, Z => n16812);
   U13891 : BUF_X1 port map( A => n15776, Z => n16803);
   U13892 : BUF_X1 port map( A => n15189, Z => n16914);
   U13893 : BUF_X1 port map( A => n15192, Z => n16905);
   U13894 : BUF_X1 port map( A => n15195, Z => n16896);
   U13895 : BUF_X1 port map( A => n15792, Z => n16767);
   U13896 : BUF_X1 port map( A => n15782, Z => n16788);
   U13897 : BUF_X1 port map( A => n15211, Z => n16860);
   U13898 : BUF_X1 port map( A => n15201, Z => n16881);
   U13899 : BUF_X1 port map( A => n15795, Z => n16758);
   U13900 : BUF_X1 port map( A => n15214, Z => n16851);
   U13901 : BUF_X1 port map( A => n17179, Z => n17172);
   U13902 : BUF_X1 port map( A => n17179, Z => n17173);
   U13903 : BUF_X1 port map( A => n17179, Z => n17174);
   U13904 : BUF_X1 port map( A => n17179, Z => n17175);
   U13905 : BUF_X1 port map( A => n17143, Z => n17136);
   U13906 : BUF_X1 port map( A => n17143, Z => n17137);
   U13907 : BUF_X1 port map( A => n17143, Z => n17138);
   U13908 : BUF_X1 port map( A => n17143, Z => n17139);
   U13909 : BUF_X1 port map( A => n17107, Z => n17100);
   U13910 : BUF_X1 port map( A => n17107, Z => n17101);
   U13911 : BUF_X1 port map( A => n17107, Z => n17102);
   U13912 : BUF_X1 port map( A => n17107, Z => n17103);
   U13913 : BUF_X1 port map( A => n17071, Z => n17064);
   U13914 : BUF_X1 port map( A => n17071, Z => n17065);
   U13915 : BUF_X1 port map( A => n17071, Z => n17066);
   U13916 : BUF_X1 port map( A => n17071, Z => n17067);
   U13917 : BUF_X1 port map( A => n17053, Z => n17046);
   U13918 : BUF_X1 port map( A => n17053, Z => n17047);
   U13919 : BUF_X1 port map( A => n17053, Z => n17048);
   U13920 : BUF_X1 port map( A => n17053, Z => n17049);
   U13921 : BUF_X1 port map( A => n17044, Z => n17037);
   U13922 : BUF_X1 port map( A => n17044, Z => n17038);
   U13923 : BUF_X1 port map( A => n17044, Z => n17039);
   U13924 : BUF_X1 port map( A => n17044, Z => n17040);
   U13925 : BUF_X1 port map( A => n17035, Z => n17028);
   U13926 : BUF_X1 port map( A => n17035, Z => n17029);
   U13927 : BUF_X1 port map( A => n17035, Z => n17030);
   U13928 : BUF_X1 port map( A => n17035, Z => n17031);
   U13929 : BUF_X1 port map( A => n17026, Z => n17019);
   U13930 : BUF_X1 port map( A => n17026, Z => n17020);
   U13931 : BUF_X1 port map( A => n17026, Z => n17021);
   U13932 : BUF_X1 port map( A => n17026, Z => n17022);
   U13933 : BUF_X1 port map( A => n17017, Z => n17010);
   U13934 : BUF_X1 port map( A => n17017, Z => n17011);
   U13935 : BUF_X1 port map( A => n17017, Z => n17012);
   U13936 : BUF_X1 port map( A => n17017, Z => n17013);
   U13937 : BUF_X1 port map( A => n17008, Z => n17001);
   U13938 : BUF_X1 port map( A => n17008, Z => n17002);
   U13939 : BUF_X1 port map( A => n17008, Z => n17003);
   U13940 : BUF_X1 port map( A => n17008, Z => n17004);
   U13941 : BUF_X1 port map( A => n16999, Z => n16992);
   U13942 : BUF_X1 port map( A => n16999, Z => n16993);
   U13943 : BUF_X1 port map( A => n16999, Z => n16994);
   U13944 : BUF_X1 port map( A => n16999, Z => n16995);
   U13945 : BUF_X1 port map( A => n16990, Z => n16983);
   U13946 : BUF_X1 port map( A => n16990, Z => n16984);
   U13947 : BUF_X1 port map( A => n16990, Z => n16985);
   U13948 : BUF_X1 port map( A => n16990, Z => n16986);
   U13949 : BUF_X1 port map( A => n16981, Z => n16974);
   U13950 : BUF_X1 port map( A => n16981, Z => n16975);
   U13951 : BUF_X1 port map( A => n16981, Z => n16976);
   U13952 : BUF_X1 port map( A => n16981, Z => n16977);
   U13953 : BUF_X1 port map( A => n16972, Z => n16965);
   U13954 : BUF_X1 port map( A => n16972, Z => n16966);
   U13955 : BUF_X1 port map( A => n16972, Z => n16967);
   U13956 : BUF_X1 port map( A => n16972, Z => n16968);
   U13957 : BUF_X1 port map( A => n16963, Z => n16956);
   U13958 : BUF_X1 port map( A => n16963, Z => n16957);
   U13959 : BUF_X1 port map( A => n16963, Z => n16958);
   U13960 : BUF_X1 port map( A => n16963, Z => n16959);
   U13961 : BUF_X1 port map( A => n16954, Z => n16947);
   U13962 : BUF_X1 port map( A => n16954, Z => n16948);
   U13963 : BUF_X1 port map( A => n16954, Z => n16949);
   U13964 : BUF_X1 port map( A => n16954, Z => n16950);
   U13965 : BUF_X1 port map( A => n16945, Z => n16938);
   U13966 : BUF_X1 port map( A => n16945, Z => n16939);
   U13967 : BUF_X1 port map( A => n16945, Z => n16940);
   U13968 : BUF_X1 port map( A => n16945, Z => n16941);
   U13969 : BUF_X1 port map( A => n16936, Z => n16929);
   U13970 : BUF_X1 port map( A => n16936, Z => n16930);
   U13971 : BUF_X1 port map( A => n16936, Z => n16931);
   U13972 : BUF_X1 port map( A => n16936, Z => n16932);
   U13973 : BUF_X1 port map( A => n17179, Z => n17176);
   U13974 : BUF_X1 port map( A => n17179, Z => n17177);
   U13975 : BUF_X1 port map( A => n17143, Z => n17140);
   U13976 : BUF_X1 port map( A => n17143, Z => n17141);
   U13977 : BUF_X1 port map( A => n17107, Z => n17104);
   U13978 : BUF_X1 port map( A => n17107, Z => n17105);
   U13979 : BUF_X1 port map( A => n17071, Z => n17068);
   U13980 : BUF_X1 port map( A => n17071, Z => n17069);
   U13981 : BUF_X1 port map( A => n17053, Z => n17050);
   U13982 : BUF_X1 port map( A => n17053, Z => n17051);
   U13983 : BUF_X1 port map( A => n17044, Z => n17041);
   U13984 : BUF_X1 port map( A => n17044, Z => n17042);
   U13985 : BUF_X1 port map( A => n17035, Z => n17032);
   U13986 : BUF_X1 port map( A => n17035, Z => n17033);
   U13987 : BUF_X1 port map( A => n17026, Z => n17023);
   U13988 : BUF_X1 port map( A => n17026, Z => n17024);
   U13989 : BUF_X1 port map( A => n17017, Z => n17014);
   U13990 : BUF_X1 port map( A => n17017, Z => n17015);
   U13991 : BUF_X1 port map( A => n17008, Z => n17005);
   U13992 : BUF_X1 port map( A => n17008, Z => n17006);
   U13993 : BUF_X1 port map( A => n16999, Z => n16996);
   U13994 : BUF_X1 port map( A => n16999, Z => n16997);
   U13995 : BUF_X1 port map( A => n16990, Z => n16987);
   U13996 : BUF_X1 port map( A => n16990, Z => n16988);
   U13997 : BUF_X1 port map( A => n16981, Z => n16978);
   U13998 : BUF_X1 port map( A => n16981, Z => n16979);
   U13999 : BUF_X1 port map( A => n16972, Z => n16969);
   U14000 : BUF_X1 port map( A => n16972, Z => n16970);
   U14001 : BUF_X1 port map( A => n16963, Z => n16960);
   U14002 : BUF_X1 port map( A => n16963, Z => n16961);
   U14003 : BUF_X1 port map( A => n16954, Z => n16951);
   U14004 : BUF_X1 port map( A => n16954, Z => n16952);
   U14005 : BUF_X1 port map( A => n16945, Z => n16942);
   U14006 : BUF_X1 port map( A => n16945, Z => n16943);
   U14007 : BUF_X1 port map( A => n16936, Z => n16933);
   U14008 : BUF_X1 port map( A => n16936, Z => n16934);
   U14009 : BUF_X1 port map( A => n17080, Z => n17073);
   U14010 : BUF_X1 port map( A => n17080, Z => n17074);
   U14011 : BUF_X1 port map( A => n17080, Z => n17075);
   U14012 : BUF_X1 port map( A => n17080, Z => n17076);
   U14013 : BUF_X1 port map( A => n17080, Z => n17077);
   U14014 : BUF_X1 port map( A => n17080, Z => n17078);
   U14015 : BUF_X1 port map( A => n17089, Z => n17082);
   U14016 : BUF_X1 port map( A => n17089, Z => n17083);
   U14017 : BUF_X1 port map( A => n17089, Z => n17084);
   U14018 : BUF_X1 port map( A => n17089, Z => n17085);
   U14019 : BUF_X1 port map( A => n17089, Z => n17086);
   U14020 : BUF_X1 port map( A => n17089, Z => n17087);
   U14021 : BUF_X1 port map( A => n17098, Z => n17091);
   U14022 : BUF_X1 port map( A => n17098, Z => n17092);
   U14023 : BUF_X1 port map( A => n17098, Z => n17093);
   U14024 : BUF_X1 port map( A => n17098, Z => n17094);
   U14025 : BUF_X1 port map( A => n17098, Z => n17095);
   U14026 : BUF_X1 port map( A => n17098, Z => n17096);
   U14027 : BUF_X1 port map( A => n17116, Z => n17109);
   U14028 : BUF_X1 port map( A => n17116, Z => n17110);
   U14029 : BUF_X1 port map( A => n17116, Z => n17111);
   U14030 : BUF_X1 port map( A => n17116, Z => n17112);
   U14031 : BUF_X1 port map( A => n17116, Z => n17113);
   U14032 : BUF_X1 port map( A => n17116, Z => n17114);
   U14033 : BUF_X1 port map( A => n17125, Z => n17118);
   U14034 : BUF_X1 port map( A => n17125, Z => n17119);
   U14035 : BUF_X1 port map( A => n17125, Z => n17120);
   U14036 : BUF_X1 port map( A => n17125, Z => n17121);
   U14037 : BUF_X1 port map( A => n17125, Z => n17122);
   U14038 : BUF_X1 port map( A => n17125, Z => n17123);
   U14039 : BUF_X1 port map( A => n17134, Z => n17127);
   U14040 : BUF_X1 port map( A => n17134, Z => n17128);
   U14041 : BUF_X1 port map( A => n17134, Z => n17129);
   U14042 : BUF_X1 port map( A => n17134, Z => n17130);
   U14043 : BUF_X1 port map( A => n17134, Z => n17131);
   U14044 : BUF_X1 port map( A => n17134, Z => n17132);
   U14045 : BUF_X1 port map( A => n17152, Z => n17145);
   U14046 : BUF_X1 port map( A => n17152, Z => n17146);
   U14047 : BUF_X1 port map( A => n17152, Z => n17147);
   U14048 : BUF_X1 port map( A => n17152, Z => n17148);
   U14049 : BUF_X1 port map( A => n17152, Z => n17149);
   U14050 : BUF_X1 port map( A => n17152, Z => n17150);
   U14051 : BUF_X1 port map( A => n17161, Z => n17154);
   U14052 : BUF_X1 port map( A => n17161, Z => n17155);
   U14053 : BUF_X1 port map( A => n17161, Z => n17156);
   U14054 : BUF_X1 port map( A => n17161, Z => n17157);
   U14055 : BUF_X1 port map( A => n17161, Z => n17158);
   U14056 : BUF_X1 port map( A => n17161, Z => n17159);
   U14057 : BUF_X1 port map( A => n17170, Z => n17163);
   U14058 : BUF_X1 port map( A => n17170, Z => n17164);
   U14059 : BUF_X1 port map( A => n17170, Z => n17165);
   U14060 : BUF_X1 port map( A => n17170, Z => n17166);
   U14061 : BUF_X1 port map( A => n17170, Z => n17167);
   U14062 : BUF_X1 port map( A => n17170, Z => n17168);
   U14063 : BUF_X1 port map( A => n17188, Z => n17181);
   U14064 : BUF_X1 port map( A => n17188, Z => n17182);
   U14065 : BUF_X1 port map( A => n17188, Z => n17183);
   U14066 : BUF_X1 port map( A => n17188, Z => n17184);
   U14067 : BUF_X1 port map( A => n17188, Z => n17185);
   U14068 : BUF_X1 port map( A => n17188, Z => n17186);
   U14069 : BUF_X1 port map( A => n17197, Z => n17190);
   U14070 : BUF_X1 port map( A => n17197, Z => n17191);
   U14071 : BUF_X1 port map( A => n17197, Z => n17192);
   U14072 : BUF_X1 port map( A => n17197, Z => n17193);
   U14073 : BUF_X1 port map( A => n17197, Z => n17194);
   U14074 : BUF_X1 port map( A => n17197, Z => n17195);
   U14075 : BUF_X1 port map( A => n17179, Z => n17178);
   U14076 : BUF_X1 port map( A => n17143, Z => n17142);
   U14077 : BUF_X1 port map( A => n17107, Z => n17106);
   U14078 : BUF_X1 port map( A => n17071, Z => n17070);
   U14079 : BUF_X1 port map( A => n17053, Z => n17052);
   U14080 : BUF_X1 port map( A => n17044, Z => n17043);
   U14081 : BUF_X1 port map( A => n17035, Z => n17034);
   U14082 : BUF_X1 port map( A => n17026, Z => n17025);
   U14083 : BUF_X1 port map( A => n17017, Z => n17016);
   U14084 : BUF_X1 port map( A => n17008, Z => n17007);
   U14085 : BUF_X1 port map( A => n16999, Z => n16998);
   U14086 : BUF_X1 port map( A => n16990, Z => n16989);
   U14087 : BUF_X1 port map( A => n16981, Z => n16980);
   U14088 : BUF_X1 port map( A => n16972, Z => n16971);
   U14089 : BUF_X1 port map( A => n16963, Z => n16962);
   U14090 : BUF_X1 port map( A => n16954, Z => n16953);
   U14091 : BUF_X1 port map( A => n16945, Z => n16944);
   U14092 : BUF_X1 port map( A => n16936, Z => n16935);
   U14093 : BUF_X1 port map( A => n17080, Z => n17079);
   U14094 : BUF_X1 port map( A => n17089, Z => n17088);
   U14095 : BUF_X1 port map( A => n17098, Z => n17097);
   U14096 : BUF_X1 port map( A => n17116, Z => n17115);
   U14097 : BUF_X1 port map( A => n17125, Z => n17124);
   U14098 : BUF_X1 port map( A => n17134, Z => n17133);
   U14099 : BUF_X1 port map( A => n17152, Z => n17151);
   U14100 : BUF_X1 port map( A => n17161, Z => n17160);
   U14101 : BUF_X1 port map( A => n17170, Z => n17169);
   U14102 : BUF_X1 port map( A => n17188, Z => n17187);
   U14103 : BUF_X1 port map( A => n17197, Z => n17196);
   U14104 : INV_X1 port map( A => n15103, ZN => n17299);
   U14105 : OAI21_X1 port map( B1 => n15135, B2 => n15136, A => n17320, ZN => 
                           n15103);
   U14106 : INV_X1 port map( A => n15159, ZN => n17062);
   U14107 : OAI21_X1 port map( B1 => n15136, B2 => n15160, A => n17318, ZN => 
                           n15159);
   U14108 : INV_X1 port map( A => n16918, ZN => n16927);
   U14109 : OAI222_X1 port map( A1 => n14820, A2 => n16815, B1 => n14757, B2 =>
                           n16812, C1 => n14597, C2 => n16809, ZN => n15918);
   U14110 : OAI222_X1 port map( A1 => n14819, A2 => n16815, B1 => n14756, B2 =>
                           n16812, C1 => n14596, C2 => n16809, ZN => n15901);
   U14111 : OAI222_X1 port map( A1 => n14818, A2 => n16815, B1 => n14755, B2 =>
                           n16812, C1 => n14595, C2 => n16809, ZN => n15884);
   U14112 : OAI222_X1 port map( A1 => n14817, A2 => n16815, B1 => n14754, B2 =>
                           n16812, C1 => n14594, C2 => n16809, ZN => n15867);
   U14113 : OAI222_X1 port map( A1 => n14816, A2 => n16815, B1 => n14753, B2 =>
                           n16812, C1 => n14593, C2 => n16809, ZN => n15850);
   U14114 : OAI222_X1 port map( A1 => n14815, A2 => n16815, B1 => n14752, B2 =>
                           n16812, C1 => n14592, C2 => n16809, ZN => n15833);
   U14115 : OAI222_X1 port map( A1 => n14814, A2 => n16815, B1 => n14751, B2 =>
                           n16812, C1 => n14591, C2 => n16809, ZN => n15816);
   U14116 : OAI222_X1 port map( A1 => n15101, A2 => n16815, B1 => n14750, B2 =>
                           n16812, C1 => n14590, C2 => n16809, ZN => n15767);
   U14117 : OAI222_X1 port map( A1 => n14820, A2 => n16908, B1 => n14757, B2 =>
                           n16905, C1 => n14597, C2 => n16902, ZN => n15337);
   U14118 : OAI222_X1 port map( A1 => n14819, A2 => n16908, B1 => n14756, B2 =>
                           n16905, C1 => n14596, C2 => n16902, ZN => n15320);
   U14119 : OAI222_X1 port map( A1 => n14818, A2 => n16908, B1 => n14755, B2 =>
                           n16905, C1 => n14595, C2 => n16902, ZN => n15303);
   U14120 : OAI222_X1 port map( A1 => n14817, A2 => n16908, B1 => n14754, B2 =>
                           n16905, C1 => n14594, C2 => n16902, ZN => n15286);
   U14121 : OAI222_X1 port map( A1 => n14816, A2 => n16908, B1 => n14753, B2 =>
                           n16905, C1 => n14593, C2 => n16902, ZN => n15269);
   U14122 : OAI222_X1 port map( A1 => n14815, A2 => n16908, B1 => n14752, B2 =>
                           n16905, C1 => n14592, C2 => n16902, ZN => n15252);
   U14123 : OAI222_X1 port map( A1 => n14814, A2 => n16908, B1 => n14751, B2 =>
                           n16905, C1 => n14591, C2 => n16902, ZN => n15235);
   U14124 : OAI222_X1 port map( A1 => n15101, A2 => n16908, B1 => n14750, B2 =>
                           n16905, C1 => n14590, C2 => n16902, ZN => n15186);
   U14125 : OAI222_X1 port map( A1 => n14844, A2 => n16813, B1 => n14781, B2 =>
                           n16810, C1 => n14621, C2 => n16807, ZN => n16326);
   U14126 : OAI222_X1 port map( A1 => n14843, A2 => n16813, B1 => n14780, B2 =>
                           n16810, C1 => n14620, C2 => n16807, ZN => n16309);
   U14127 : OAI222_X1 port map( A1 => n14842, A2 => n16813, B1 => n14779, B2 =>
                           n16810, C1 => n14619, C2 => n16807, ZN => n16292);
   U14128 : OAI222_X1 port map( A1 => n14841, A2 => n16813, B1 => n14778, B2 =>
                           n16810, C1 => n14618, C2 => n16807, ZN => n16275);
   U14129 : OAI222_X1 port map( A1 => n14840, A2 => n16813, B1 => n14777, B2 =>
                           n16810, C1 => n14617, C2 => n16807, ZN => n16258);
   U14130 : OAI222_X1 port map( A1 => n14839, A2 => n16813, B1 => n14776, B2 =>
                           n16810, C1 => n14616, C2 => n16807, ZN => n16241);
   U14131 : OAI222_X1 port map( A1 => n14838, A2 => n16813, B1 => n14775, B2 =>
                           n16810, C1 => n14615, C2 => n16807, ZN => n16224);
   U14132 : OAI222_X1 port map( A1 => n14837, A2 => n16813, B1 => n14774, B2 =>
                           n16810, C1 => n14614, C2 => n16807, ZN => n16207);
   U14133 : OAI222_X1 port map( A1 => n14836, A2 => n16813, B1 => n14773, B2 =>
                           n16810, C1 => n14613, C2 => n16807, ZN => n16190);
   U14134 : OAI222_X1 port map( A1 => n14835, A2 => n16813, B1 => n14772, B2 =>
                           n16810, C1 => n14612, C2 => n16807, ZN => n16173);
   U14135 : OAI222_X1 port map( A1 => n14834, A2 => n16813, B1 => n14771, B2 =>
                           n16810, C1 => n14611, C2 => n16807, ZN => n16156);
   U14136 : OAI222_X1 port map( A1 => n14833, A2 => n16813, B1 => n14770, B2 =>
                           n16810, C1 => n14610, C2 => n16807, ZN => n16139);
   U14137 : OAI222_X1 port map( A1 => n14832, A2 => n16814, B1 => n14769, B2 =>
                           n16811, C1 => n14609, C2 => n16808, ZN => n16122);
   U14138 : OAI222_X1 port map( A1 => n14831, A2 => n16814, B1 => n14768, B2 =>
                           n16811, C1 => n14608, C2 => n16808, ZN => n16105);
   U14139 : OAI222_X1 port map( A1 => n14830, A2 => n16814, B1 => n14767, B2 =>
                           n16811, C1 => n14607, C2 => n16808, ZN => n16088);
   U14140 : OAI222_X1 port map( A1 => n14829, A2 => n16814, B1 => n14766, B2 =>
                           n16811, C1 => n14606, C2 => n16808, ZN => n16071);
   U14141 : OAI222_X1 port map( A1 => n14828, A2 => n16814, B1 => n14765, B2 =>
                           n16811, C1 => n14605, C2 => n16808, ZN => n16054);
   U14142 : OAI222_X1 port map( A1 => n14827, A2 => n16814, B1 => n14764, B2 =>
                           n16811, C1 => n14604, C2 => n16808, ZN => n16037);
   U14143 : OAI222_X1 port map( A1 => n14826, A2 => n16814, B1 => n14763, B2 =>
                           n16811, C1 => n14603, C2 => n16808, ZN => n16020);
   U14144 : OAI222_X1 port map( A1 => n14825, A2 => n16814, B1 => n14762, B2 =>
                           n16811, C1 => n14602, C2 => n16808, ZN => n16003);
   U14145 : OAI222_X1 port map( A1 => n14824, A2 => n16814, B1 => n14761, B2 =>
                           n16811, C1 => n14601, C2 => n16808, ZN => n15986);
   U14146 : OAI222_X1 port map( A1 => n14823, A2 => n16814, B1 => n14760, B2 =>
                           n16811, C1 => n14600, C2 => n16808, ZN => n15969);
   U14147 : OAI222_X1 port map( A1 => n14822, A2 => n16814, B1 => n14759, B2 =>
                           n16811, C1 => n14599, C2 => n16808, ZN => n15952);
   U14148 : OAI222_X1 port map( A1 => n14821, A2 => n16814, B1 => n14758, B2 =>
                           n16811, C1 => n14598, C2 => n16808, ZN => n15935);
   U14149 : OAI222_X1 port map( A1 => n14844, A2 => n16906, B1 => n14781, B2 =>
                           n16903, C1 => n14621, C2 => n16900, ZN => n15745);
   U14150 : OAI222_X1 port map( A1 => n14843, A2 => n16906, B1 => n14780, B2 =>
                           n16903, C1 => n14620, C2 => n16900, ZN => n15728);
   U14151 : OAI222_X1 port map( A1 => n14842, A2 => n16906, B1 => n14779, B2 =>
                           n16903, C1 => n14619, C2 => n16900, ZN => n15711);
   U14152 : OAI222_X1 port map( A1 => n14841, A2 => n16906, B1 => n14778, B2 =>
                           n16903, C1 => n14618, C2 => n16900, ZN => n15694);
   U14153 : OAI222_X1 port map( A1 => n14840, A2 => n16906, B1 => n14777, B2 =>
                           n16903, C1 => n14617, C2 => n16900, ZN => n15677);
   U14154 : OAI222_X1 port map( A1 => n14839, A2 => n16906, B1 => n14776, B2 =>
                           n16903, C1 => n14616, C2 => n16900, ZN => n15660);
   U14155 : OAI222_X1 port map( A1 => n14838, A2 => n16906, B1 => n14775, B2 =>
                           n16903, C1 => n14615, C2 => n16900, ZN => n15643);
   U14156 : OAI222_X1 port map( A1 => n14837, A2 => n16906, B1 => n14774, B2 =>
                           n16903, C1 => n14614, C2 => n16900, ZN => n15626);
   U14157 : OAI222_X1 port map( A1 => n14836, A2 => n16906, B1 => n14773, B2 =>
                           n16903, C1 => n14613, C2 => n16900, ZN => n15609);
   U14158 : OAI222_X1 port map( A1 => n14835, A2 => n16906, B1 => n14772, B2 =>
                           n16903, C1 => n14612, C2 => n16900, ZN => n15592);
   U14159 : OAI222_X1 port map( A1 => n14834, A2 => n16906, B1 => n14771, B2 =>
                           n16903, C1 => n14611, C2 => n16900, ZN => n15575);
   U14160 : OAI222_X1 port map( A1 => n14833, A2 => n16906, B1 => n14770, B2 =>
                           n16903, C1 => n14610, C2 => n16900, ZN => n15558);
   U14161 : OAI222_X1 port map( A1 => n14832, A2 => n16907, B1 => n14769, B2 =>
                           n16904, C1 => n14609, C2 => n16901, ZN => n15541);
   U14162 : OAI222_X1 port map( A1 => n14831, A2 => n16907, B1 => n14768, B2 =>
                           n16904, C1 => n14608, C2 => n16901, ZN => n15524);
   U14163 : OAI222_X1 port map( A1 => n14830, A2 => n16907, B1 => n14767, B2 =>
                           n16904, C1 => n14607, C2 => n16901, ZN => n15507);
   U14164 : OAI222_X1 port map( A1 => n14829, A2 => n16907, B1 => n14766, B2 =>
                           n16904, C1 => n14606, C2 => n16901, ZN => n15490);
   U14165 : OAI222_X1 port map( A1 => n14828, A2 => n16907, B1 => n14765, B2 =>
                           n16904, C1 => n14605, C2 => n16901, ZN => n15473);
   U14166 : OAI222_X1 port map( A1 => n14827, A2 => n16907, B1 => n14764, B2 =>
                           n16904, C1 => n14604, C2 => n16901, ZN => n15456);
   U14167 : OAI222_X1 port map( A1 => n14826, A2 => n16907, B1 => n14763, B2 =>
                           n16904, C1 => n14603, C2 => n16901, ZN => n15439);
   U14168 : OAI222_X1 port map( A1 => n14825, A2 => n16907, B1 => n14762, B2 =>
                           n16904, C1 => n14602, C2 => n16901, ZN => n15422);
   U14169 : OAI222_X1 port map( A1 => n14824, A2 => n16907, B1 => n14761, B2 =>
                           n16904, C1 => n14601, C2 => n16901, ZN => n15405);
   U14170 : OAI222_X1 port map( A1 => n14823, A2 => n16907, B1 => n14760, B2 =>
                           n16904, C1 => n14600, C2 => n16901, ZN => n15388);
   U14171 : OAI222_X1 port map( A1 => n14822, A2 => n16907, B1 => n14759, B2 =>
                           n16904, C1 => n14599, C2 => n16901, ZN => n15371);
   U14172 : OAI222_X1 port map( A1 => n14821, A2 => n16907, B1 => n14758, B2 =>
                           n16904, C1 => n14598, C2 => n16901, ZN => n15354);
   U14173 : OAI22_X1 port map( A1 => n17079, A2 => n17301, B1 => n15157, B2 => 
                           n15101, ZN => n1915);
   U14174 : OAI22_X1 port map( A1 => n17077, A2 => n17271, B1 => n15157, B2 => 
                           n14820, ZN => n1908);
   U14175 : OAI22_X1 port map( A1 => n17078, A2 => n17274, B1 => n15157, B2 => 
                           n14819, ZN => n1909);
   U14176 : OAI22_X1 port map( A1 => n17078, A2 => n17277, B1 => n15157, B2 => 
                           n14818, ZN => n1910);
   U14177 : OAI22_X1 port map( A1 => n17078, A2 => n17280, B1 => n15157, B2 => 
                           n14817, ZN => n1911);
   U14178 : OAI22_X1 port map( A1 => n17078, A2 => n17283, B1 => n15157, B2 => 
                           n14816, ZN => n1912);
   U14179 : OAI22_X1 port map( A1 => n17078, A2 => n17286, B1 => n15157, B2 => 
                           n14815, ZN => n1913);
   U14180 : OAI22_X1 port map( A1 => n17079, A2 => n17289, B1 => n15157, B2 => 
                           n14814, ZN => n1914);
   U14181 : OAI22_X1 port map( A1 => n17086, A2 => n17271, B1 => n15156, B2 => 
                           n14789, ZN => n1940);
   U14182 : OAI22_X1 port map( A1 => n17087, A2 => n17274, B1 => n15156, B2 => 
                           n14788, ZN => n1941);
   U14183 : OAI22_X1 port map( A1 => n17087, A2 => n17277, B1 => n15156, B2 => 
                           n14787, ZN => n1942);
   U14184 : OAI22_X1 port map( A1 => n17087, A2 => n17280, B1 => n15156, B2 => 
                           n14786, ZN => n1943);
   U14185 : OAI22_X1 port map( A1 => n17087, A2 => n17283, B1 => n15156, B2 => 
                           n14785, ZN => n1944);
   U14186 : OAI22_X1 port map( A1 => n17087, A2 => n17286, B1 => n15156, B2 => 
                           n14784, ZN => n1945);
   U14187 : OAI22_X1 port map( A1 => n17088, A2 => n17289, B1 => n15156, B2 => 
                           n14783, ZN => n1946);
   U14188 : OAI22_X1 port map( A1 => n17088, A2 => n17301, B1 => n15156, B2 => 
                           n14782, ZN => n1947);
   U14189 : OAI22_X1 port map( A1 => n17095, A2 => n17271, B1 => n15154, B2 => 
                           n14757, ZN => n1972);
   U14190 : OAI22_X1 port map( A1 => n17096, A2 => n17274, B1 => n15154, B2 => 
                           n14756, ZN => n1973);
   U14191 : OAI22_X1 port map( A1 => n17096, A2 => n17277, B1 => n15154, B2 => 
                           n14755, ZN => n1974);
   U14192 : OAI22_X1 port map( A1 => n17096, A2 => n17280, B1 => n15154, B2 => 
                           n14754, ZN => n1975);
   U14193 : OAI22_X1 port map( A1 => n17096, A2 => n17283, B1 => n15154, B2 => 
                           n14753, ZN => n1976);
   U14194 : OAI22_X1 port map( A1 => n17096, A2 => n17286, B1 => n15154, B2 => 
                           n14752, ZN => n1977);
   U14195 : OAI22_X1 port map( A1 => n17097, A2 => n17289, B1 => n15154, B2 => 
                           n14751, ZN => n1978);
   U14196 : OAI22_X1 port map( A1 => n17097, A2 => n17301, B1 => n15154, B2 => 
                           n14750, ZN => n1979);
   U14197 : OAI22_X1 port map( A1 => n17122, A2 => n17270, B1 => n15151, B2 => 
                           n14693, ZN => n2068);
   U14198 : OAI22_X1 port map( A1 => n17123, A2 => n17273, B1 => n15151, B2 => 
                           n14692, ZN => n2069);
   U14199 : OAI22_X1 port map( A1 => n17123, A2 => n17276, B1 => n15151, B2 => 
                           n14691, ZN => n2070);
   U14200 : OAI22_X1 port map( A1 => n17123, A2 => n17279, B1 => n15151, B2 => 
                           n14690, ZN => n2071);
   U14201 : OAI22_X1 port map( A1 => n17123, A2 => n17282, B1 => n15151, B2 => 
                           n14689, ZN => n2072);
   U14202 : OAI22_X1 port map( A1 => n17123, A2 => n17285, B1 => n15151, B2 => 
                           n14688, ZN => n2073);
   U14203 : OAI22_X1 port map( A1 => n17124, A2 => n17288, B1 => n15151, B2 => 
                           n14687, ZN => n2074);
   U14204 : OAI22_X1 port map( A1 => n17124, A2 => n17300, B1 => n15151, B2 => 
                           n14686, ZN => n2075);
   U14205 : OAI22_X1 port map( A1 => n17149, A2 => n17270, B1 => n15147, B2 => 
                           n14629, ZN => n2164);
   U14206 : OAI22_X1 port map( A1 => n17150, A2 => n17273, B1 => n15147, B2 => 
                           n14628, ZN => n2165);
   U14207 : OAI22_X1 port map( A1 => n17150, A2 => n17276, B1 => n15147, B2 => 
                           n14627, ZN => n2166);
   U14208 : OAI22_X1 port map( A1 => n17150, A2 => n17279, B1 => n15147, B2 => 
                           n14626, ZN => n2167);
   U14209 : OAI22_X1 port map( A1 => n17150, A2 => n17282, B1 => n15147, B2 => 
                           n14625, ZN => n2168);
   U14210 : OAI22_X1 port map( A1 => n17150, A2 => n17285, B1 => n15147, B2 => 
                           n14624, ZN => n2169);
   U14211 : OAI22_X1 port map( A1 => n17151, A2 => n17288, B1 => n15147, B2 => 
                           n14623, ZN => n2170);
   U14212 : OAI22_X1 port map( A1 => n17151, A2 => n17300, B1 => n15147, B2 => 
                           n14622, ZN => n2171);
   U14213 : OAI22_X1 port map( A1 => n17158, A2 => n17270, B1 => n15146, B2 => 
                           n14597, ZN => n2196);
   U14214 : OAI22_X1 port map( A1 => n17159, A2 => n17273, B1 => n15146, B2 => 
                           n14596, ZN => n2197);
   U14215 : OAI22_X1 port map( A1 => n17159, A2 => n17276, B1 => n15146, B2 => 
                           n14595, ZN => n2198);
   U14216 : OAI22_X1 port map( A1 => n17159, A2 => n17279, B1 => n15146, B2 => 
                           n14594, ZN => n2199);
   U14217 : OAI22_X1 port map( A1 => n17159, A2 => n17282, B1 => n15146, B2 => 
                           n14593, ZN => n2200);
   U14218 : OAI22_X1 port map( A1 => n17159, A2 => n17285, B1 => n15146, B2 => 
                           n14592, ZN => n2201);
   U14219 : OAI22_X1 port map( A1 => n17160, A2 => n17288, B1 => n15146, B2 => 
                           n14591, ZN => n2202);
   U14220 : OAI22_X1 port map( A1 => n17160, A2 => n17300, B1 => n15146, B2 => 
                           n14590, ZN => n2203);
   U14221 : OAI22_X1 port map( A1 => n17167, A2 => n17270, B1 => n15144, B2 => 
                           n14565, ZN => n2228);
   U14222 : OAI22_X1 port map( A1 => n17168, A2 => n17273, B1 => n15144, B2 => 
                           n14564, ZN => n2229);
   U14223 : OAI22_X1 port map( A1 => n17168, A2 => n17276, B1 => n15144, B2 => 
                           n14563, ZN => n2230);
   U14224 : OAI22_X1 port map( A1 => n17168, A2 => n17279, B1 => n15144, B2 => 
                           n14562, ZN => n2231);
   U14225 : OAI22_X1 port map( A1 => n17168, A2 => n17282, B1 => n15144, B2 => 
                           n14561, ZN => n2232);
   U14226 : OAI22_X1 port map( A1 => n17168, A2 => n17285, B1 => n15144, B2 => 
                           n14560, ZN => n2233);
   U14227 : OAI22_X1 port map( A1 => n17169, A2 => n17288, B1 => n15144, B2 => 
                           n14559, ZN => n2234);
   U14228 : OAI22_X1 port map( A1 => n17169, A2 => n17300, B1 => n15144, B2 => 
                           n14558, ZN => n2235);
   U14229 : OAI22_X1 port map( A1 => n17073, A2 => n17199, B1 => n17072, B2 => 
                           n14844, ZN => n1884);
   U14230 : OAI22_X1 port map( A1 => n17073, A2 => n17202, B1 => n17072, B2 => 
                           n14843, ZN => n1885);
   U14231 : OAI22_X1 port map( A1 => n17073, A2 => n17205, B1 => n17072, B2 => 
                           n14842, ZN => n1886);
   U14232 : OAI22_X1 port map( A1 => n17073, A2 => n17208, B1 => n17072, B2 => 
                           n14841, ZN => n1887);
   U14233 : OAI22_X1 port map( A1 => n17073, A2 => n17211, B1 => n17072, B2 => 
                           n14840, ZN => n1888);
   U14234 : OAI22_X1 port map( A1 => n17074, A2 => n17214, B1 => n17072, B2 => 
                           n14839, ZN => n1889);
   U14235 : OAI22_X1 port map( A1 => n17074, A2 => n17217, B1 => n17072, B2 => 
                           n14838, ZN => n1890);
   U14236 : OAI22_X1 port map( A1 => n17074, A2 => n17220, B1 => n17072, B2 => 
                           n14837, ZN => n1891);
   U14237 : OAI22_X1 port map( A1 => n17074, A2 => n17223, B1 => n17072, B2 => 
                           n14836, ZN => n1892);
   U14238 : OAI22_X1 port map( A1 => n17074, A2 => n17226, B1 => n17072, B2 => 
                           n14835, ZN => n1893);
   U14239 : OAI22_X1 port map( A1 => n17075, A2 => n17229, B1 => n17072, B2 => 
                           n14834, ZN => n1894);
   U14240 : OAI22_X1 port map( A1 => n17075, A2 => n17232, B1 => n17072, B2 => 
                           n14833, ZN => n1895);
   U14241 : OAI22_X1 port map( A1 => n17075, A2 => n17235, B1 => n15157, B2 => 
                           n14832, ZN => n1896);
   U14242 : OAI22_X1 port map( A1 => n17075, A2 => n17238, B1 => n15157, B2 => 
                           n14831, ZN => n1897);
   U14243 : OAI22_X1 port map( A1 => n17075, A2 => n17241, B1 => n15157, B2 => 
                           n14830, ZN => n1898);
   U14244 : OAI22_X1 port map( A1 => n17076, A2 => n17244, B1 => n17072, B2 => 
                           n14829, ZN => n1899);
   U14245 : OAI22_X1 port map( A1 => n17076, A2 => n17247, B1 => n17072, B2 => 
                           n14828, ZN => n1900);
   U14246 : OAI22_X1 port map( A1 => n17076, A2 => n17250, B1 => n17072, B2 => 
                           n14827, ZN => n1901);
   U14247 : OAI22_X1 port map( A1 => n17076, A2 => n17253, B1 => n17072, B2 => 
                           n14826, ZN => n1902);
   U14248 : OAI22_X1 port map( A1 => n17076, A2 => n17256, B1 => n17072, B2 => 
                           n14825, ZN => n1903);
   U14249 : OAI22_X1 port map( A1 => n17077, A2 => n17259, B1 => n17072, B2 => 
                           n14824, ZN => n1904);
   U14250 : OAI22_X1 port map( A1 => n17077, A2 => n17262, B1 => n17072, B2 => 
                           n14823, ZN => n1905);
   U14251 : OAI22_X1 port map( A1 => n17077, A2 => n17265, B1 => n17072, B2 => 
                           n14822, ZN => n1906);
   U14252 : OAI22_X1 port map( A1 => n17077, A2 => n17268, B1 => n17072, B2 => 
                           n14821, ZN => n1907);
   U14253 : OAI22_X1 port map( A1 => n17082, A2 => n17199, B1 => n17081, B2 => 
                           n14813, ZN => n1916);
   U14254 : OAI22_X1 port map( A1 => n17082, A2 => n17202, B1 => n17081, B2 => 
                           n14812, ZN => n1917);
   U14255 : OAI22_X1 port map( A1 => n17082, A2 => n17205, B1 => n17081, B2 => 
                           n14811, ZN => n1918);
   U14256 : OAI22_X1 port map( A1 => n17082, A2 => n17208, B1 => n17081, B2 => 
                           n14810, ZN => n1919);
   U14257 : OAI22_X1 port map( A1 => n17082, A2 => n17211, B1 => n17081, B2 => 
                           n14809, ZN => n1920);
   U14258 : OAI22_X1 port map( A1 => n17083, A2 => n17214, B1 => n17081, B2 => 
                           n14808, ZN => n1921);
   U14259 : OAI22_X1 port map( A1 => n17083, A2 => n17217, B1 => n17081, B2 => 
                           n14807, ZN => n1922);
   U14260 : OAI22_X1 port map( A1 => n17083, A2 => n17220, B1 => n17081, B2 => 
                           n14806, ZN => n1923);
   U14261 : OAI22_X1 port map( A1 => n17083, A2 => n17223, B1 => n17081, B2 => 
                           n14805, ZN => n1924);
   U14262 : OAI22_X1 port map( A1 => n17083, A2 => n17226, B1 => n17081, B2 => 
                           n14804, ZN => n1925);
   U14263 : OAI22_X1 port map( A1 => n17084, A2 => n17229, B1 => n17081, B2 => 
                           n14803, ZN => n1926);
   U14264 : OAI22_X1 port map( A1 => n17084, A2 => n17232, B1 => n17081, B2 => 
                           n14802, ZN => n1927);
   U14265 : OAI22_X1 port map( A1 => n17084, A2 => n17235, B1 => n15156, B2 => 
                           n14801, ZN => n1928);
   U14266 : OAI22_X1 port map( A1 => n17084, A2 => n17238, B1 => n15156, B2 => 
                           n14800, ZN => n1929);
   U14267 : OAI22_X1 port map( A1 => n17084, A2 => n17241, B1 => n15156, B2 => 
                           n14799, ZN => n1930);
   U14268 : OAI22_X1 port map( A1 => n17085, A2 => n17244, B1 => n17081, B2 => 
                           n14798, ZN => n1931);
   U14269 : OAI22_X1 port map( A1 => n17085, A2 => n17247, B1 => n17081, B2 => 
                           n14797, ZN => n1932);
   U14270 : OAI22_X1 port map( A1 => n17085, A2 => n17250, B1 => n17081, B2 => 
                           n14796, ZN => n1933);
   U14271 : OAI22_X1 port map( A1 => n17085, A2 => n17253, B1 => n17081, B2 => 
                           n14795, ZN => n1934);
   U14272 : OAI22_X1 port map( A1 => n17085, A2 => n17256, B1 => n17081, B2 => 
                           n14794, ZN => n1935);
   U14273 : OAI22_X1 port map( A1 => n17086, A2 => n17259, B1 => n17081, B2 => 
                           n14793, ZN => n1936);
   U14274 : OAI22_X1 port map( A1 => n17086, A2 => n17262, B1 => n17081, B2 => 
                           n14792, ZN => n1937);
   U14275 : OAI22_X1 port map( A1 => n17086, A2 => n17265, B1 => n17081, B2 => 
                           n14791, ZN => n1938);
   U14276 : OAI22_X1 port map( A1 => n17086, A2 => n17268, B1 => n17081, B2 => 
                           n14790, ZN => n1939);
   U14277 : OAI22_X1 port map( A1 => n17091, A2 => n17199, B1 => n17090, B2 => 
                           n14781, ZN => n1948);
   U14278 : OAI22_X1 port map( A1 => n17091, A2 => n17202, B1 => n17090, B2 => 
                           n14780, ZN => n1949);
   U14279 : OAI22_X1 port map( A1 => n17091, A2 => n17205, B1 => n17090, B2 => 
                           n14779, ZN => n1950);
   U14280 : OAI22_X1 port map( A1 => n17091, A2 => n17208, B1 => n17090, B2 => 
                           n14778, ZN => n1951);
   U14281 : OAI22_X1 port map( A1 => n17091, A2 => n17211, B1 => n17090, B2 => 
                           n14777, ZN => n1952);
   U14282 : OAI22_X1 port map( A1 => n17092, A2 => n17214, B1 => n17090, B2 => 
                           n14776, ZN => n1953);
   U14283 : OAI22_X1 port map( A1 => n17092, A2 => n17217, B1 => n17090, B2 => 
                           n14775, ZN => n1954);
   U14284 : OAI22_X1 port map( A1 => n17092, A2 => n17220, B1 => n17090, B2 => 
                           n14774, ZN => n1955);
   U14285 : OAI22_X1 port map( A1 => n17092, A2 => n17223, B1 => n17090, B2 => 
                           n14773, ZN => n1956);
   U14286 : OAI22_X1 port map( A1 => n17092, A2 => n17226, B1 => n17090, B2 => 
                           n14772, ZN => n1957);
   U14287 : OAI22_X1 port map( A1 => n17093, A2 => n17229, B1 => n17090, B2 => 
                           n14771, ZN => n1958);
   U14288 : OAI22_X1 port map( A1 => n17093, A2 => n17232, B1 => n17090, B2 => 
                           n14770, ZN => n1959);
   U14289 : OAI22_X1 port map( A1 => n17093, A2 => n17235, B1 => n15154, B2 => 
                           n14769, ZN => n1960);
   U14290 : OAI22_X1 port map( A1 => n17093, A2 => n17238, B1 => n15154, B2 => 
                           n14768, ZN => n1961);
   U14291 : OAI22_X1 port map( A1 => n17093, A2 => n17241, B1 => n15154, B2 => 
                           n14767, ZN => n1962);
   U14292 : OAI22_X1 port map( A1 => n17094, A2 => n17244, B1 => n17090, B2 => 
                           n14766, ZN => n1963);
   U14293 : OAI22_X1 port map( A1 => n17094, A2 => n17247, B1 => n17090, B2 => 
                           n14765, ZN => n1964);
   U14294 : OAI22_X1 port map( A1 => n17094, A2 => n17250, B1 => n17090, B2 => 
                           n14764, ZN => n1965);
   U14295 : OAI22_X1 port map( A1 => n17094, A2 => n17253, B1 => n17090, B2 => 
                           n14763, ZN => n1966);
   U14296 : OAI22_X1 port map( A1 => n17094, A2 => n17256, B1 => n17090, B2 => 
                           n14762, ZN => n1967);
   U14297 : OAI22_X1 port map( A1 => n17095, A2 => n17259, B1 => n17090, B2 => 
                           n14761, ZN => n1968);
   U14298 : OAI22_X1 port map( A1 => n17095, A2 => n17262, B1 => n17090, B2 => 
                           n14760, ZN => n1969);
   U14299 : OAI22_X1 port map( A1 => n17095, A2 => n17265, B1 => n17090, B2 => 
                           n14759, ZN => n1970);
   U14300 : OAI22_X1 port map( A1 => n17095, A2 => n17268, B1 => n17090, B2 => 
                           n14758, ZN => n1971);
   U14301 : OAI22_X1 port map( A1 => n17118, A2 => n17198, B1 => n17117, B2 => 
                           n14717, ZN => n2044);
   U14302 : OAI22_X1 port map( A1 => n17118, A2 => n17201, B1 => n17117, B2 => 
                           n14716, ZN => n2045);
   U14303 : OAI22_X1 port map( A1 => n17118, A2 => n17204, B1 => n17117, B2 => 
                           n14715, ZN => n2046);
   U14304 : OAI22_X1 port map( A1 => n17118, A2 => n17207, B1 => n17117, B2 => 
                           n14714, ZN => n2047);
   U14305 : OAI22_X1 port map( A1 => n17118, A2 => n17210, B1 => n17117, B2 => 
                           n14713, ZN => n2048);
   U14306 : OAI22_X1 port map( A1 => n17119, A2 => n17213, B1 => n17117, B2 => 
                           n14712, ZN => n2049);
   U14307 : OAI22_X1 port map( A1 => n17119, A2 => n17216, B1 => n17117, B2 => 
                           n14711, ZN => n2050);
   U14308 : OAI22_X1 port map( A1 => n17119, A2 => n17219, B1 => n17117, B2 => 
                           n14710, ZN => n2051);
   U14309 : OAI22_X1 port map( A1 => n17119, A2 => n17222, B1 => n17117, B2 => 
                           n14709, ZN => n2052);
   U14310 : OAI22_X1 port map( A1 => n17119, A2 => n17225, B1 => n17117, B2 => 
                           n14708, ZN => n2053);
   U14311 : OAI22_X1 port map( A1 => n17120, A2 => n17228, B1 => n17117, B2 => 
                           n14707, ZN => n2054);
   U14312 : OAI22_X1 port map( A1 => n17120, A2 => n17231, B1 => n17117, B2 => 
                           n14706, ZN => n2055);
   U14313 : OAI22_X1 port map( A1 => n17120, A2 => n17234, B1 => n15151, B2 => 
                           n14705, ZN => n2056);
   U14314 : OAI22_X1 port map( A1 => n17120, A2 => n17237, B1 => n15151, B2 => 
                           n14704, ZN => n2057);
   U14315 : OAI22_X1 port map( A1 => n17120, A2 => n17240, B1 => n15151, B2 => 
                           n14703, ZN => n2058);
   U14316 : OAI22_X1 port map( A1 => n17121, A2 => n17243, B1 => n17117, B2 => 
                           n14702, ZN => n2059);
   U14317 : OAI22_X1 port map( A1 => n17121, A2 => n17246, B1 => n17117, B2 => 
                           n14701, ZN => n2060);
   U14318 : OAI22_X1 port map( A1 => n17121, A2 => n17249, B1 => n17117, B2 => 
                           n14700, ZN => n2061);
   U14319 : OAI22_X1 port map( A1 => n17121, A2 => n17252, B1 => n17117, B2 => 
                           n14699, ZN => n2062);
   U14320 : OAI22_X1 port map( A1 => n17121, A2 => n17255, B1 => n17117, B2 => 
                           n14698, ZN => n2063);
   U14321 : OAI22_X1 port map( A1 => n17122, A2 => n17258, B1 => n17117, B2 => 
                           n14697, ZN => n2064);
   U14322 : OAI22_X1 port map( A1 => n17122, A2 => n17261, B1 => n17117, B2 => 
                           n14696, ZN => n2065);
   U14323 : OAI22_X1 port map( A1 => n17122, A2 => n17264, B1 => n17117, B2 => 
                           n14695, ZN => n2066);
   U14324 : OAI22_X1 port map( A1 => n17122, A2 => n17267, B1 => n17117, B2 => 
                           n14694, ZN => n2067);
   U14325 : OAI22_X1 port map( A1 => n17145, A2 => n17198, B1 => n17144, B2 => 
                           n14653, ZN => n2140);
   U14326 : OAI22_X1 port map( A1 => n17145, A2 => n17201, B1 => n17144, B2 => 
                           n14652, ZN => n2141);
   U14327 : OAI22_X1 port map( A1 => n17145, A2 => n17204, B1 => n17144, B2 => 
                           n14651, ZN => n2142);
   U14328 : OAI22_X1 port map( A1 => n17145, A2 => n17207, B1 => n17144, B2 => 
                           n14650, ZN => n2143);
   U14329 : OAI22_X1 port map( A1 => n17145, A2 => n17210, B1 => n17144, B2 => 
                           n14649, ZN => n2144);
   U14330 : OAI22_X1 port map( A1 => n17146, A2 => n17213, B1 => n17144, B2 => 
                           n14648, ZN => n2145);
   U14331 : OAI22_X1 port map( A1 => n17146, A2 => n17216, B1 => n17144, B2 => 
                           n14647, ZN => n2146);
   U14332 : OAI22_X1 port map( A1 => n17146, A2 => n17219, B1 => n17144, B2 => 
                           n14646, ZN => n2147);
   U14333 : OAI22_X1 port map( A1 => n17146, A2 => n17222, B1 => n17144, B2 => 
                           n14645, ZN => n2148);
   U14334 : OAI22_X1 port map( A1 => n17146, A2 => n17225, B1 => n17144, B2 => 
                           n14644, ZN => n2149);
   U14335 : OAI22_X1 port map( A1 => n17147, A2 => n17228, B1 => n17144, B2 => 
                           n14643, ZN => n2150);
   U14336 : OAI22_X1 port map( A1 => n17147, A2 => n17231, B1 => n17144, B2 => 
                           n14642, ZN => n2151);
   U14337 : OAI22_X1 port map( A1 => n17147, A2 => n17234, B1 => n15147, B2 => 
                           n14641, ZN => n2152);
   U14338 : OAI22_X1 port map( A1 => n17147, A2 => n17237, B1 => n15147, B2 => 
                           n14640, ZN => n2153);
   U14339 : OAI22_X1 port map( A1 => n17147, A2 => n17240, B1 => n15147, B2 => 
                           n14639, ZN => n2154);
   U14340 : OAI22_X1 port map( A1 => n17148, A2 => n17243, B1 => n17144, B2 => 
                           n14638, ZN => n2155);
   U14341 : OAI22_X1 port map( A1 => n17148, A2 => n17246, B1 => n17144, B2 => 
                           n14637, ZN => n2156);
   U14342 : OAI22_X1 port map( A1 => n17148, A2 => n17249, B1 => n17144, B2 => 
                           n14636, ZN => n2157);
   U14343 : OAI22_X1 port map( A1 => n17148, A2 => n17252, B1 => n17144, B2 => 
                           n14635, ZN => n2158);
   U14344 : OAI22_X1 port map( A1 => n17148, A2 => n17255, B1 => n17144, B2 => 
                           n14634, ZN => n2159);
   U14345 : OAI22_X1 port map( A1 => n17149, A2 => n17258, B1 => n17144, B2 => 
                           n14633, ZN => n2160);
   U14346 : OAI22_X1 port map( A1 => n17149, A2 => n17261, B1 => n17144, B2 => 
                           n14632, ZN => n2161);
   U14347 : OAI22_X1 port map( A1 => n17149, A2 => n17264, B1 => n17144, B2 => 
                           n14631, ZN => n2162);
   U14348 : OAI22_X1 port map( A1 => n17149, A2 => n17267, B1 => n17144, B2 => 
                           n14630, ZN => n2163);
   U14349 : OAI22_X1 port map( A1 => n17154, A2 => n17198, B1 => n17153, B2 => 
                           n14621, ZN => n2172);
   U14350 : OAI22_X1 port map( A1 => n17154, A2 => n17201, B1 => n17153, B2 => 
                           n14620, ZN => n2173);
   U14351 : OAI22_X1 port map( A1 => n17154, A2 => n17204, B1 => n17153, B2 => 
                           n14619, ZN => n2174);
   U14352 : OAI22_X1 port map( A1 => n17154, A2 => n17207, B1 => n17153, B2 => 
                           n14618, ZN => n2175);
   U14353 : OAI22_X1 port map( A1 => n17154, A2 => n17210, B1 => n17153, B2 => 
                           n14617, ZN => n2176);
   U14354 : OAI22_X1 port map( A1 => n17155, A2 => n17213, B1 => n17153, B2 => 
                           n14616, ZN => n2177);
   U14355 : OAI22_X1 port map( A1 => n17155, A2 => n17216, B1 => n17153, B2 => 
                           n14615, ZN => n2178);
   U14356 : OAI22_X1 port map( A1 => n17155, A2 => n17219, B1 => n17153, B2 => 
                           n14614, ZN => n2179);
   U14357 : OAI22_X1 port map( A1 => n17155, A2 => n17222, B1 => n17153, B2 => 
                           n14613, ZN => n2180);
   U14358 : OAI22_X1 port map( A1 => n17155, A2 => n17225, B1 => n17153, B2 => 
                           n14612, ZN => n2181);
   U14359 : OAI22_X1 port map( A1 => n17156, A2 => n17228, B1 => n17153, B2 => 
                           n14611, ZN => n2182);
   U14360 : OAI22_X1 port map( A1 => n17156, A2 => n17231, B1 => n17153, B2 => 
                           n14610, ZN => n2183);
   U14361 : OAI22_X1 port map( A1 => n17156, A2 => n17234, B1 => n15146, B2 => 
                           n14609, ZN => n2184);
   U14362 : OAI22_X1 port map( A1 => n17156, A2 => n17237, B1 => n15146, B2 => 
                           n14608, ZN => n2185);
   U14363 : OAI22_X1 port map( A1 => n17156, A2 => n17240, B1 => n15146, B2 => 
                           n14607, ZN => n2186);
   U14364 : OAI22_X1 port map( A1 => n17157, A2 => n17243, B1 => n17153, B2 => 
                           n14606, ZN => n2187);
   U14365 : OAI22_X1 port map( A1 => n17157, A2 => n17246, B1 => n17153, B2 => 
                           n14605, ZN => n2188);
   U14366 : OAI22_X1 port map( A1 => n17157, A2 => n17249, B1 => n17153, B2 => 
                           n14604, ZN => n2189);
   U14367 : OAI22_X1 port map( A1 => n17157, A2 => n17252, B1 => n17153, B2 => 
                           n14603, ZN => n2190);
   U14368 : OAI22_X1 port map( A1 => n17157, A2 => n17255, B1 => n17153, B2 => 
                           n14602, ZN => n2191);
   U14369 : OAI22_X1 port map( A1 => n17158, A2 => n17258, B1 => n17153, B2 => 
                           n14601, ZN => n2192);
   U14370 : OAI22_X1 port map( A1 => n17158, A2 => n17261, B1 => n17153, B2 => 
                           n14600, ZN => n2193);
   U14371 : OAI22_X1 port map( A1 => n17158, A2 => n17264, B1 => n17153, B2 => 
                           n14599, ZN => n2194);
   U14372 : OAI22_X1 port map( A1 => n17158, A2 => n17267, B1 => n17153, B2 => 
                           n14598, ZN => n2195);
   U14373 : OAI22_X1 port map( A1 => n17163, A2 => n17198, B1 => n17162, B2 => 
                           n14589, ZN => n2204);
   U14374 : OAI22_X1 port map( A1 => n17163, A2 => n17201, B1 => n17162, B2 => 
                           n14588, ZN => n2205);
   U14375 : OAI22_X1 port map( A1 => n17163, A2 => n17204, B1 => n17162, B2 => 
                           n14587, ZN => n2206);
   U14376 : OAI22_X1 port map( A1 => n17163, A2 => n17207, B1 => n17162, B2 => 
                           n14586, ZN => n2207);
   U14377 : OAI22_X1 port map( A1 => n17163, A2 => n17210, B1 => n17162, B2 => 
                           n14585, ZN => n2208);
   U14378 : OAI22_X1 port map( A1 => n17164, A2 => n17213, B1 => n17162, B2 => 
                           n14584, ZN => n2209);
   U14379 : OAI22_X1 port map( A1 => n17164, A2 => n17216, B1 => n17162, B2 => 
                           n14583, ZN => n2210);
   U14380 : OAI22_X1 port map( A1 => n17164, A2 => n17219, B1 => n17162, B2 => 
                           n14582, ZN => n2211);
   U14381 : OAI22_X1 port map( A1 => n17164, A2 => n17222, B1 => n17162, B2 => 
                           n14581, ZN => n2212);
   U14382 : OAI22_X1 port map( A1 => n17164, A2 => n17225, B1 => n17162, B2 => 
                           n14580, ZN => n2213);
   U14383 : OAI22_X1 port map( A1 => n17165, A2 => n17228, B1 => n17162, B2 => 
                           n14579, ZN => n2214);
   U14384 : OAI22_X1 port map( A1 => n17165, A2 => n17231, B1 => n17162, B2 => 
                           n14578, ZN => n2215);
   U14385 : OAI22_X1 port map( A1 => n17165, A2 => n17234, B1 => n15144, B2 => 
                           n14577, ZN => n2216);
   U14386 : OAI22_X1 port map( A1 => n17165, A2 => n17237, B1 => n15144, B2 => 
                           n14576, ZN => n2217);
   U14387 : OAI22_X1 port map( A1 => n17165, A2 => n17240, B1 => n15144, B2 => 
                           n14575, ZN => n2218);
   U14388 : OAI22_X1 port map( A1 => n17166, A2 => n17243, B1 => n17162, B2 => 
                           n14574, ZN => n2219);
   U14389 : OAI22_X1 port map( A1 => n17166, A2 => n17246, B1 => n17162, B2 => 
                           n14573, ZN => n2220);
   U14390 : OAI22_X1 port map( A1 => n17166, A2 => n17249, B1 => n17162, B2 => 
                           n14572, ZN => n2221);
   U14391 : OAI22_X1 port map( A1 => n17166, A2 => n17252, B1 => n17162, B2 => 
                           n14571, ZN => n2222);
   U14392 : OAI22_X1 port map( A1 => n17166, A2 => n17255, B1 => n17162, B2 => 
                           n14570, ZN => n2223);
   U14393 : OAI22_X1 port map( A1 => n17167, A2 => n17258, B1 => n17162, B2 => 
                           n14569, ZN => n2224);
   U14394 : OAI22_X1 port map( A1 => n17167, A2 => n17261, B1 => n17162, B2 => 
                           n14568, ZN => n2225);
   U14395 : OAI22_X1 port map( A1 => n17167, A2 => n17264, B1 => n17162, B2 => 
                           n14567, ZN => n2226);
   U14396 : OAI22_X1 port map( A1 => n17167, A2 => n17267, B1 => n17162, B2 => 
                           n14566, ZN => n2227);
   U14397 : INV_X1 port map( A => n16726, ZN => n16754);
   U14398 : INV_X1 port map( A => n16727, ZN => n16847);
   U14399 : INV_X1 port map( A => n16728, ZN => n16740);
   U14400 : INV_X1 port map( A => n16728, ZN => n16741);
   U14401 : INV_X1 port map( A => n16729, ZN => n16833);
   U14402 : INV_X1 port map( A => n16729, ZN => n16834);
   U14403 : INV_X1 port map( A => n16730, ZN => n16738);
   U14404 : INV_X1 port map( A => n16731, ZN => n16831);
   U14405 : NAND2_X1 port map( A1 => n14446, A2 => n14447, ZN => n15136);
   U14406 : BUF_X1 port map( A => n15807, Z => n16735);
   U14407 : BUF_X1 port map( A => n15807, Z => n16736);
   U14408 : BUF_X1 port map( A => n15226, Z => n16828);
   U14409 : BUF_X1 port map( A => n15226, Z => n16829);
   U14410 : BUF_X1 port map( A => n15808, Z => n16732);
   U14411 : BUF_X1 port map( A => n15808, Z => n16733);
   U14412 : BUF_X1 port map( A => n15227, Z => n16825);
   U14413 : BUF_X1 port map( A => n15227, Z => n16826);
   U14414 : NAND2_X1 port map( A1 => n16331, A2 => n16730, ZN => n15778);
   U14415 : NAND2_X1 port map( A1 => n15750, A2 => n16731, ZN => n15197);
   U14416 : BUF_X1 port map( A => n15807, Z => n16737);
   U14417 : BUF_X1 port map( A => n15226, Z => n16830);
   U14418 : BUF_X1 port map( A => n14442, Z => n17319);
   U14419 : BUF_X1 port map( A => n14442, Z => n17318);
   U14420 : INV_X1 port map( A => n16726, ZN => n16755);
   U14421 : INV_X1 port map( A => n16727, ZN => n16848);
   U14422 : BUF_X1 port map( A => n15808, Z => n16734);
   U14423 : BUF_X1 port map( A => n15227, Z => n16827);
   U14424 : BUF_X1 port map( A => n14442, Z => n17316);
   U14425 : BUF_X1 port map( A => n14442, Z => n17315);
   U14426 : BUF_X1 port map( A => n15134, Z => n17199);
   U14427 : BUF_X1 port map( A => n15133, Z => n17202);
   U14428 : BUF_X1 port map( A => n15132, Z => n17205);
   U14429 : BUF_X1 port map( A => n15131, Z => n17208);
   U14430 : BUF_X1 port map( A => n15130, Z => n17211);
   U14431 : BUF_X1 port map( A => n15129, Z => n17214);
   U14432 : BUF_X1 port map( A => n15128, Z => n17217);
   U14433 : BUF_X1 port map( A => n15127, Z => n17220);
   U14434 : BUF_X1 port map( A => n15126, Z => n17223);
   U14435 : BUF_X1 port map( A => n15125, Z => n17226);
   U14436 : BUF_X1 port map( A => n15124, Z => n17229);
   U14437 : BUF_X1 port map( A => n15123, Z => n17232);
   U14438 : BUF_X1 port map( A => n15122, Z => n17235);
   U14439 : BUF_X1 port map( A => n15121, Z => n17238);
   U14440 : BUF_X1 port map( A => n15120, Z => n17241);
   U14441 : BUF_X1 port map( A => n15119, Z => n17244);
   U14442 : BUF_X1 port map( A => n15118, Z => n17247);
   U14443 : BUF_X1 port map( A => n15117, Z => n17250);
   U14444 : BUF_X1 port map( A => n15116, Z => n17253);
   U14445 : BUF_X1 port map( A => n15115, Z => n17256);
   U14446 : BUF_X1 port map( A => n15114, Z => n17259);
   U14447 : BUF_X1 port map( A => n15113, Z => n17262);
   U14448 : BUF_X1 port map( A => n15112, Z => n17265);
   U14449 : BUF_X1 port map( A => n15111, Z => n17268);
   U14450 : BUF_X1 port map( A => n15110, Z => n17271);
   U14451 : BUF_X1 port map( A => n15109, Z => n17274);
   U14452 : BUF_X1 port map( A => n15108, Z => n17277);
   U14453 : BUF_X1 port map( A => n15107, Z => n17280);
   U14454 : BUF_X1 port map( A => n15106, Z => n17283);
   U14455 : BUF_X1 port map( A => n15105, Z => n17286);
   U14456 : BUF_X1 port map( A => n15104, Z => n17289);
   U14457 : BUF_X1 port map( A => n15102, Z => n17301);
   U14458 : BUF_X1 port map( A => n15134, Z => n17198);
   U14459 : BUF_X1 port map( A => n15133, Z => n17201);
   U14460 : BUF_X1 port map( A => n15132, Z => n17204);
   U14461 : BUF_X1 port map( A => n15131, Z => n17207);
   U14462 : BUF_X1 port map( A => n15130, Z => n17210);
   U14463 : BUF_X1 port map( A => n15129, Z => n17213);
   U14464 : BUF_X1 port map( A => n15128, Z => n17216);
   U14465 : BUF_X1 port map( A => n15127, Z => n17219);
   U14466 : BUF_X1 port map( A => n15126, Z => n17222);
   U14467 : BUF_X1 port map( A => n15125, Z => n17225);
   U14468 : BUF_X1 port map( A => n15124, Z => n17228);
   U14469 : BUF_X1 port map( A => n15123, Z => n17231);
   U14470 : BUF_X1 port map( A => n15122, Z => n17234);
   U14471 : BUF_X1 port map( A => n15121, Z => n17237);
   U14472 : BUF_X1 port map( A => n15120, Z => n17240);
   U14473 : BUF_X1 port map( A => n15119, Z => n17243);
   U14474 : BUF_X1 port map( A => n15118, Z => n17246);
   U14475 : BUF_X1 port map( A => n15117, Z => n17249);
   U14476 : BUF_X1 port map( A => n15116, Z => n17252);
   U14477 : BUF_X1 port map( A => n15115, Z => n17255);
   U14478 : BUF_X1 port map( A => n15114, Z => n17258);
   U14479 : BUF_X1 port map( A => n15113, Z => n17261);
   U14480 : BUF_X1 port map( A => n15112, Z => n17264);
   U14481 : BUF_X1 port map( A => n15111, Z => n17267);
   U14482 : BUF_X1 port map( A => n15110, Z => n17270);
   U14483 : BUF_X1 port map( A => n15109, Z => n17273);
   U14484 : BUF_X1 port map( A => n15108, Z => n17276);
   U14485 : BUF_X1 port map( A => n15107, Z => n17279);
   U14486 : BUF_X1 port map( A => n15106, Z => n17282);
   U14487 : BUF_X1 port map( A => n15105, Z => n17285);
   U14488 : BUF_X1 port map( A => n15104, Z => n17288);
   U14489 : BUF_X1 port map( A => n15102, Z => n17300);
   U14490 : BUF_X1 port map( A => n14442, Z => n17317);
   U14491 : BUF_X1 port map( A => n15802, Z => n16745);
   U14492 : BUF_X1 port map( A => n15802, Z => n16746);
   U14493 : BUF_X1 port map( A => n15221, Z => n16838);
   U14494 : BUF_X1 port map( A => n15221, Z => n16839);
   U14495 : BUF_X1 port map( A => n15803, Z => n16742);
   U14496 : BUF_X1 port map( A => n15803, Z => n16743);
   U14497 : BUF_X1 port map( A => n15222, Z => n16835);
   U14498 : BUF_X1 port map( A => n15222, Z => n16836);
   U14499 : BUF_X1 port map( A => n15801, Z => n16748);
   U14500 : BUF_X1 port map( A => n15801, Z => n16749);
   U14501 : BUF_X1 port map( A => n15220, Z => n16841);
   U14502 : BUF_X1 port map( A => n15220, Z => n16842);
   U14503 : BUF_X1 port map( A => n15134, Z => n17200);
   U14504 : BUF_X1 port map( A => n15133, Z => n17203);
   U14505 : BUF_X1 port map( A => n15132, Z => n17206);
   U14506 : BUF_X1 port map( A => n15131, Z => n17209);
   U14507 : BUF_X1 port map( A => n15130, Z => n17212);
   U14508 : BUF_X1 port map( A => n15129, Z => n17215);
   U14509 : BUF_X1 port map( A => n15128, Z => n17218);
   U14510 : BUF_X1 port map( A => n15127, Z => n17221);
   U14511 : BUF_X1 port map( A => n15126, Z => n17224);
   U14512 : BUF_X1 port map( A => n15125, Z => n17227);
   U14513 : BUF_X1 port map( A => n15124, Z => n17230);
   U14514 : BUF_X1 port map( A => n15123, Z => n17233);
   U14515 : BUF_X1 port map( A => n15122, Z => n17236);
   U14516 : BUF_X1 port map( A => n15121, Z => n17239);
   U14517 : BUF_X1 port map( A => n15120, Z => n17242);
   U14518 : BUF_X1 port map( A => n15119, Z => n17245);
   U14519 : BUF_X1 port map( A => n15118, Z => n17248);
   U14520 : BUF_X1 port map( A => n15117, Z => n17251);
   U14521 : BUF_X1 port map( A => n15116, Z => n17254);
   U14522 : BUF_X1 port map( A => n15115, Z => n17257);
   U14523 : BUF_X1 port map( A => n15114, Z => n17260);
   U14524 : BUF_X1 port map( A => n15113, Z => n17263);
   U14525 : BUF_X1 port map( A => n15112, Z => n17266);
   U14526 : BUF_X1 port map( A => n15111, Z => n17269);
   U14527 : BUF_X1 port map( A => n15110, Z => n17272);
   U14528 : BUF_X1 port map( A => n15109, Z => n17275);
   U14529 : BUF_X1 port map( A => n15108, Z => n17278);
   U14530 : BUF_X1 port map( A => n15107, Z => n17281);
   U14531 : BUF_X1 port map( A => n15106, Z => n17284);
   U14532 : BUF_X1 port map( A => n15105, Z => n17287);
   U14533 : BUF_X1 port map( A => n15104, Z => n17290);
   U14534 : BUF_X1 port map( A => n15102, Z => n17302);
   U14535 : BUF_X1 port map( A => n15801, Z => n16750);
   U14536 : BUF_X1 port map( A => n15220, Z => n16843);
   U14537 : BUF_X1 port map( A => n15802, Z => n16747);
   U14538 : BUF_X1 port map( A => n15221, Z => n16840);
   U14539 : BUF_X1 port map( A => n15803, Z => n16744);
   U14540 : BUF_X1 port map( A => n15222, Z => n16837);
   U14541 : NAND2_X1 port map( A1 => n16328, A2 => n16331, ZN => n15789);
   U14542 : NAND2_X1 port map( A1 => n16335, A2 => n16331, ZN => n15787);
   U14543 : NAND2_X1 port map( A1 => n16744, A2 => n16331, ZN => n15769);
   U14544 : NAND2_X1 port map( A1 => n16747, A2 => n16331, ZN => n15772);
   U14545 : NAND2_X1 port map( A1 => n16728, A2 => n16331, ZN => n15775);
   U14546 : NAND2_X1 port map( A1 => n15747, A2 => n15750, ZN => n15208);
   U14547 : NAND2_X1 port map( A1 => n15754, A2 => n15750, ZN => n15206);
   U14548 : NAND2_X1 port map( A1 => n16837, A2 => n15750, ZN => n15188);
   U14549 : NAND2_X1 port map( A1 => n16840, A2 => n15750, ZN => n15191);
   U14550 : NAND2_X1 port map( A1 => n16729, A2 => n15750, ZN => n15194);
   U14551 : NAND2_X1 port map( A1 => n16328, A2 => n16330, ZN => n15788);
   U14552 : NAND2_X1 port map( A1 => n16744, A2 => n16330, ZN => n15770);
   U14553 : NAND2_X1 port map( A1 => n16747, A2 => n16330, ZN => n15773);
   U14554 : NAND2_X1 port map( A1 => n16728, A2 => n16330, ZN => n15776);
   U14555 : NAND2_X1 port map( A1 => n15747, A2 => n15749, ZN => n15207);
   U14556 : NAND2_X1 port map( A1 => n16837, A2 => n15749, ZN => n15189);
   U14557 : NAND2_X1 port map( A1 => n16840, A2 => n15749, ZN => n15192);
   U14558 : NAND2_X1 port map( A1 => n16729, A2 => n15749, ZN => n15195);
   U14559 : NAND2_X1 port map( A1 => n16328, A2 => n16329, ZN => n15771);
   U14560 : NAND2_X1 port map( A1 => n15747, A2 => n15748, ZN => n15190);
   U14561 : NAND2_X1 port map( A1 => n16737, A2 => n16329, ZN => n15786);
   U14562 : NAND2_X1 port map( A1 => n16830, A2 => n15748, ZN => n15205);
   U14563 : INV_X1 port map( A => n16328, ZN => n14458);
   U14564 : INV_X1 port map( A => n15747, ZN => n14451);
   U14565 : AND2_X1 port map( A1 => n16330, A2 => n16730, ZN => n15782);
   U14566 : AND2_X1 port map( A1 => n15749, A2 => n16731, ZN => n15201);
   U14567 : AND2_X1 port map( A1 => n16734, A2 => n16331, ZN => n15797);
   U14568 : AND2_X1 port map( A1 => n16737, A2 => n16331, ZN => n15794);
   U14569 : AND2_X1 port map( A1 => n16827, A2 => n15750, ZN => n15216);
   U14570 : AND2_X1 port map( A1 => n16830, A2 => n15750, ZN => n15213);
   U14571 : NAND2_X1 port map( A1 => n16728, A2 => n16329, ZN => n15779);
   U14572 : NAND2_X1 port map( A1 => n16744, A2 => n16329, ZN => n15774);
   U14573 : NAND2_X1 port map( A1 => n16747, A2 => n16329, ZN => n15777);
   U14574 : NAND2_X1 port map( A1 => n16729, A2 => n15748, ZN => n15198);
   U14575 : NAND2_X1 port map( A1 => n16837, A2 => n15748, ZN => n15193);
   U14576 : NAND2_X1 port map( A1 => n16840, A2 => n15748, ZN => n15196);
   U14577 : INV_X1 port map( A => n16335, ZN => n14457);
   U14578 : INV_X1 port map( A => n15754, ZN => n14450);
   U14579 : AND2_X1 port map( A1 => n16335, A2 => n16330, ZN => n15792);
   U14580 : AND2_X1 port map( A1 => n15754, A2 => n15749, ZN => n15211);
   U14581 : AND2_X1 port map( A1 => n16737, A2 => n16330, ZN => n15783);
   U14582 : AND2_X1 port map( A1 => n16734, A2 => n16330, ZN => n15793);
   U14583 : AND2_X1 port map( A1 => n16830, A2 => n15749, ZN => n15202);
   U14584 : AND2_X1 port map( A1 => n16827, A2 => n15749, ZN => n15212);
   U14585 : AND2_X1 port map( A1 => n16335, A2 => n16329, ZN => n15791);
   U14586 : AND2_X1 port map( A1 => n15754, A2 => n15748, ZN => n15210);
   U14587 : AND2_X1 port map( A1 => n16734, A2 => n16329, ZN => n15795);
   U14588 : AND2_X1 port map( A1 => n16827, A2 => n15748, ZN => n15214);
   U14589 : AND2_X1 port map( A1 => n16730, A2 => n16329, ZN => n15781);
   U14590 : AND2_X1 port map( A1 => n16731, A2 => n15748, ZN => n15200);
   U14591 : BUF_X1 port map( A => n15179, Z => n16918);
   U14592 : OAI21_X1 port map( B1 => n15142, B2 => n15176, A => n17319, ZN => 
                           n15179);
   U14593 : INV_X1 port map( A => n15141, ZN => n17179);
   U14594 : OAI21_X1 port map( B1 => n15135, B2 => n15142, A => n17319, ZN => 
                           n15141);
   U14595 : INV_X1 port map( A => n15139, ZN => n17188);
   U14596 : OAI21_X1 port map( B1 => n15135, B2 => n15140, A => n17319, ZN => 
                           n15139);
   U14597 : INV_X1 port map( A => n15137, ZN => n17197);
   U14598 : OAI21_X1 port map( B1 => n15135, B2 => n15138, A => n17320, ZN => 
                           n15137);
   U14599 : INV_X1 port map( A => n15148, ZN => n17143);
   U14600 : OAI21_X1 port map( B1 => n15142, B2 => n15145, A => n17319, ZN => 
                           n15148);
   U14601 : INV_X1 port map( A => n15153, ZN => n17107);
   U14602 : OAI21_X1 port map( B1 => n15142, B2 => n15150, A => n17319, ZN => 
                           n15153);
   U14603 : INV_X1 port map( A => n15158, ZN => n17071);
   U14604 : OAI21_X1 port map( B1 => n15142, B2 => n15155, A => n17318, ZN => 
                           n15158);
   U14605 : INV_X1 port map( A => n15161, ZN => n17053);
   U14606 : OAI21_X1 port map( B1 => n15138, B2 => n15160, A => n17318, ZN => 
                           n15161);
   U14607 : INV_X1 port map( A => n15162, ZN => n17044);
   U14608 : OAI21_X1 port map( B1 => n15140, B2 => n15160, A => n17318, ZN => 
                           n15162);
   U14609 : INV_X1 port map( A => n15163, ZN => n17035);
   U14610 : OAI21_X1 port map( B1 => n15142, B2 => n15160, A => n17318, ZN => 
                           n15163);
   U14611 : INV_X1 port map( A => n15165, ZN => n17026);
   U14612 : OAI21_X1 port map( B1 => n15136, B2 => n15166, A => n17318, ZN => 
                           n15165);
   U14613 : INV_X1 port map( A => n15167, ZN => n17017);
   U14614 : OAI21_X1 port map( B1 => n15138, B2 => n15166, A => n17318, ZN => 
                           n15167);
   U14615 : INV_X1 port map( A => n15168, ZN => n17008);
   U14616 : OAI21_X1 port map( B1 => n15140, B2 => n15166, A => n17318, ZN => 
                           n15168);
   U14617 : INV_X1 port map( A => n15169, ZN => n16999);
   U14618 : OAI21_X1 port map( B1 => n15142, B2 => n15166, A => n17318, ZN => 
                           n15169);
   U14619 : INV_X1 port map( A => n15170, ZN => n16990);
   U14620 : OAI21_X1 port map( B1 => n15136, B2 => n15171, A => n17318, ZN => 
                           n15170);
   U14621 : INV_X1 port map( A => n15172, ZN => n16981);
   U14622 : OAI21_X1 port map( B1 => n15138, B2 => n15171, A => n17318, ZN => 
                           n15172);
   U14623 : INV_X1 port map( A => n15173, ZN => n16972);
   U14624 : OAI21_X1 port map( B1 => n15140, B2 => n15171, A => n17317, ZN => 
                           n15173);
   U14625 : INV_X1 port map( A => n15174, ZN => n16963);
   U14626 : OAI21_X1 port map( B1 => n15142, B2 => n15171, A => n17318, ZN => 
                           n15174);
   U14627 : INV_X1 port map( A => n15175, ZN => n16954);
   U14628 : OAI21_X1 port map( B1 => n15136, B2 => n15176, A => n17317, ZN => 
                           n15175);
   U14629 : INV_X1 port map( A => n15177, ZN => n16945);
   U14630 : OAI21_X1 port map( B1 => n15138, B2 => n15176, A => n17317, ZN => 
                           n15177);
   U14631 : INV_X1 port map( A => n15178, ZN => n16936);
   U14632 : OAI21_X1 port map( B1 => n15140, B2 => n15176, A => n17317, ZN => 
                           n15178);
   U14633 : INV_X1 port map( A => n15157, ZN => n17080);
   U14634 : OAI21_X1 port map( B1 => n15140, B2 => n15155, A => n17318, ZN => 
                           n15157);
   U14635 : INV_X1 port map( A => n15156, ZN => n17089);
   U14636 : OAI21_X1 port map( B1 => n15138, B2 => n15155, A => n17319, ZN => 
                           n15156);
   U14637 : INV_X1 port map( A => n15154, ZN => n17098);
   U14638 : OAI21_X1 port map( B1 => n15136, B2 => n15155, A => n17319, ZN => 
                           n15154);
   U14639 : INV_X1 port map( A => n15152, ZN => n17116);
   U14640 : OAI21_X1 port map( B1 => n15140, B2 => n15150, A => n17319, ZN => 
                           n15152);
   U14641 : INV_X1 port map( A => n15151, ZN => n17125);
   U14642 : OAI21_X1 port map( B1 => n15138, B2 => n15150, A => n17319, ZN => 
                           n15151);
   U14643 : INV_X1 port map( A => n15149, ZN => n17134);
   U14644 : OAI21_X1 port map( B1 => n15136, B2 => n15150, A => n17319, ZN => 
                           n15149);
   U14645 : INV_X1 port map( A => n15147, ZN => n17152);
   U14646 : OAI21_X1 port map( B1 => n15140, B2 => n15145, A => n17319, ZN => 
                           n15147);
   U14647 : INV_X1 port map( A => n15146, ZN => n17161);
   U14648 : OAI21_X1 port map( B1 => n15138, B2 => n15145, A => n17319, ZN => 
                           n15146);
   U14649 : INV_X1 port map( A => n15144, ZN => n17170);
   U14650 : OAI21_X1 port map( B1 => n15136, B2 => n15145, A => n17319, ZN => 
                           n15144);
   U14651 : OAI222_X1 port map( A1 => n14653, A2 => n16822, B1 => n14589, B2 =>
                           n16819, C1 => n13561, C2 => n16816, ZN => n16327);
   U14652 : OAI222_X1 port map( A1 => n14652, A2 => n16822, B1 => n14588, B2 =>
                           n16819, C1 => n13560, C2 => n16816, ZN => n16310);
   U14653 : OAI222_X1 port map( A1 => n14651, A2 => n16822, B1 => n14587, B2 =>
                           n16819, C1 => n13559, C2 => n16816, ZN => n16293);
   U14654 : OAI222_X1 port map( A1 => n14650, A2 => n16822, B1 => n14586, B2 =>
                           n16819, C1 => n13558, C2 => n16816, ZN => n16276);
   U14655 : OAI222_X1 port map( A1 => n14649, A2 => n16822, B1 => n14585, B2 =>
                           n16819, C1 => n13557, C2 => n16816, ZN => n16259);
   U14656 : OAI222_X1 port map( A1 => n14648, A2 => n16822, B1 => n14584, B2 =>
                           n16819, C1 => n13556, C2 => n16816, ZN => n16242);
   U14657 : OAI222_X1 port map( A1 => n14647, A2 => n16822, B1 => n14583, B2 =>
                           n16819, C1 => n13555, C2 => n16816, ZN => n16225);
   U14658 : OAI222_X1 port map( A1 => n14646, A2 => n16822, B1 => n14582, B2 =>
                           n16819, C1 => n13554, C2 => n16816, ZN => n16208);
   U14659 : OAI222_X1 port map( A1 => n14645, A2 => n16822, B1 => n14581, B2 =>
                           n16819, C1 => n13553, C2 => n16816, ZN => n16191);
   U14660 : OAI222_X1 port map( A1 => n14644, A2 => n16822, B1 => n14580, B2 =>
                           n16819, C1 => n13552, C2 => n16816, ZN => n16174);
   U14661 : OAI222_X1 port map( A1 => n14643, A2 => n16822, B1 => n14579, B2 =>
                           n16819, C1 => n13551, C2 => n16816, ZN => n16157);
   U14662 : OAI222_X1 port map( A1 => n14642, A2 => n16822, B1 => n14578, B2 =>
                           n16819, C1 => n13550, C2 => n16816, ZN => n16140);
   U14663 : OAI222_X1 port map( A1 => n14641, A2 => n16823, B1 => n14577, B2 =>
                           n16820, C1 => n13549, C2 => n16817, ZN => n16123);
   U14664 : OAI222_X1 port map( A1 => n14640, A2 => n16823, B1 => n14576, B2 =>
                           n16820, C1 => n13548, C2 => n16817, ZN => n16106);
   U14665 : OAI222_X1 port map( A1 => n14639, A2 => n16823, B1 => n14575, B2 =>
                           n16820, C1 => n13547, C2 => n16817, ZN => n16089);
   U14666 : OAI222_X1 port map( A1 => n14638, A2 => n16823, B1 => n14574, B2 =>
                           n16820, C1 => n13546, C2 => n16817, ZN => n16072);
   U14667 : OAI222_X1 port map( A1 => n14637, A2 => n16823, B1 => n14573, B2 =>
                           n16820, C1 => n13545, C2 => n16817, ZN => n16055);
   U14668 : OAI222_X1 port map( A1 => n14636, A2 => n16823, B1 => n14572, B2 =>
                           n16820, C1 => n13544, C2 => n16817, ZN => n16038);
   U14669 : OAI222_X1 port map( A1 => n14635, A2 => n16823, B1 => n14571, B2 =>
                           n16820, C1 => n13543, C2 => n16817, ZN => n16021);
   U14670 : OAI222_X1 port map( A1 => n14634, A2 => n16823, B1 => n14570, B2 =>
                           n16820, C1 => n13542, C2 => n16817, ZN => n16004);
   U14671 : OAI222_X1 port map( A1 => n14633, A2 => n16823, B1 => n14569, B2 =>
                           n16820, C1 => n13541, C2 => n16817, ZN => n15987);
   U14672 : OAI222_X1 port map( A1 => n14632, A2 => n16823, B1 => n14568, B2 =>
                           n16820, C1 => n13540, C2 => n16817, ZN => n15970);
   U14673 : OAI222_X1 port map( A1 => n14631, A2 => n16823, B1 => n14567, B2 =>
                           n16820, C1 => n13539, C2 => n16817, ZN => n15953);
   U14674 : OAI222_X1 port map( A1 => n14630, A2 => n16823, B1 => n14566, B2 =>
                           n16820, C1 => n13538, C2 => n16817, ZN => n15936);
   U14675 : OAI222_X1 port map( A1 => n14629, A2 => n16824, B1 => n14565, B2 =>
                           n16821, C1 => n13537, C2 => n16818, ZN => n15919);
   U14676 : OAI222_X1 port map( A1 => n14628, A2 => n16824, B1 => n14564, B2 =>
                           n16821, C1 => n13536, C2 => n16818, ZN => n15902);
   U14677 : OAI222_X1 port map( A1 => n14627, A2 => n16824, B1 => n14563, B2 =>
                           n16821, C1 => n13535, C2 => n16818, ZN => n15885);
   U14678 : OAI222_X1 port map( A1 => n14626, A2 => n16824, B1 => n14562, B2 =>
                           n16821, C1 => n13534, C2 => n16818, ZN => n15868);
   U14679 : OAI222_X1 port map( A1 => n14625, A2 => n16824, B1 => n14561, B2 =>
                           n16821, C1 => n13533, C2 => n16818, ZN => n15851);
   U14680 : OAI222_X1 port map( A1 => n14624, A2 => n16824, B1 => n14560, B2 =>
                           n16821, C1 => n13532, C2 => n16818, ZN => n15834);
   U14681 : OAI222_X1 port map( A1 => n14623, A2 => n16824, B1 => n14559, B2 =>
                           n16821, C1 => n13531, C2 => n16818, ZN => n15817);
   U14682 : OAI222_X1 port map( A1 => n14622, A2 => n16824, B1 => n14558, B2 =>
                           n16821, C1 => n13530, C2 => n16818, ZN => n15768);
   U14683 : OAI222_X1 port map( A1 => n14653, A2 => n16915, B1 => n14589, B2 =>
                           n16912, C1 => n13561, C2 => n16909, ZN => n15746);
   U14684 : OAI222_X1 port map( A1 => n14652, A2 => n16915, B1 => n14588, B2 =>
                           n16912, C1 => n13560, C2 => n16909, ZN => n15729);
   U14685 : OAI222_X1 port map( A1 => n14651, A2 => n16915, B1 => n14587, B2 =>
                           n16912, C1 => n13559, C2 => n16909, ZN => n15712);
   U14686 : OAI222_X1 port map( A1 => n14650, A2 => n16915, B1 => n14586, B2 =>
                           n16912, C1 => n13558, C2 => n16909, ZN => n15695);
   U14687 : OAI222_X1 port map( A1 => n14649, A2 => n16915, B1 => n14585, B2 =>
                           n16912, C1 => n13557, C2 => n16909, ZN => n15678);
   U14688 : OAI222_X1 port map( A1 => n14648, A2 => n16915, B1 => n14584, B2 =>
                           n16912, C1 => n13556, C2 => n16909, ZN => n15661);
   U14689 : OAI222_X1 port map( A1 => n14647, A2 => n16915, B1 => n14583, B2 =>
                           n16912, C1 => n13555, C2 => n16909, ZN => n15644);
   U14690 : OAI222_X1 port map( A1 => n14646, A2 => n16915, B1 => n14582, B2 =>
                           n16912, C1 => n13554, C2 => n16909, ZN => n15627);
   U14691 : OAI222_X1 port map( A1 => n14645, A2 => n16915, B1 => n14581, B2 =>
                           n16912, C1 => n13553, C2 => n16909, ZN => n15610);
   U14692 : OAI222_X1 port map( A1 => n14644, A2 => n16915, B1 => n14580, B2 =>
                           n16912, C1 => n13552, C2 => n16909, ZN => n15593);
   U14693 : OAI222_X1 port map( A1 => n14643, A2 => n16915, B1 => n14579, B2 =>
                           n16912, C1 => n13551, C2 => n16909, ZN => n15576);
   U14694 : OAI222_X1 port map( A1 => n14642, A2 => n16915, B1 => n14578, B2 =>
                           n16912, C1 => n13550, C2 => n16909, ZN => n15559);
   U14695 : OAI222_X1 port map( A1 => n14641, A2 => n16916, B1 => n14577, B2 =>
                           n16913, C1 => n13549, C2 => n16910, ZN => n15542);
   U14696 : OAI222_X1 port map( A1 => n14640, A2 => n16916, B1 => n14576, B2 =>
                           n16913, C1 => n13548, C2 => n16910, ZN => n15525);
   U14697 : OAI222_X1 port map( A1 => n14639, A2 => n16916, B1 => n14575, B2 =>
                           n16913, C1 => n13547, C2 => n16910, ZN => n15508);
   U14698 : OAI222_X1 port map( A1 => n14638, A2 => n16916, B1 => n14574, B2 =>
                           n16913, C1 => n13546, C2 => n16910, ZN => n15491);
   U14699 : OAI222_X1 port map( A1 => n14637, A2 => n16916, B1 => n14573, B2 =>
                           n16913, C1 => n13545, C2 => n16910, ZN => n15474);
   U14700 : OAI222_X1 port map( A1 => n14636, A2 => n16916, B1 => n14572, B2 =>
                           n16913, C1 => n13544, C2 => n16910, ZN => n15457);
   U14701 : OAI222_X1 port map( A1 => n14635, A2 => n16916, B1 => n14571, B2 =>
                           n16913, C1 => n13543, C2 => n16910, ZN => n15440);
   U14702 : OAI222_X1 port map( A1 => n14634, A2 => n16916, B1 => n14570, B2 =>
                           n16913, C1 => n13542, C2 => n16910, ZN => n15423);
   U14703 : OAI222_X1 port map( A1 => n14633, A2 => n16916, B1 => n14569, B2 =>
                           n16913, C1 => n13541, C2 => n16910, ZN => n15406);
   U14704 : OAI222_X1 port map( A1 => n14632, A2 => n16916, B1 => n14568, B2 =>
                           n16913, C1 => n13540, C2 => n16910, ZN => n15389);
   U14705 : OAI222_X1 port map( A1 => n14631, A2 => n16916, B1 => n14567, B2 =>
                           n16913, C1 => n13539, C2 => n16910, ZN => n15372);
   U14706 : OAI222_X1 port map( A1 => n14630, A2 => n16916, B1 => n14566, B2 =>
                           n16913, C1 => n13538, C2 => n16910, ZN => n15355);
   U14707 : OAI222_X1 port map( A1 => n14629, A2 => n16917, B1 => n14565, B2 =>
                           n16914, C1 => n13537, C2 => n16911, ZN => n15338);
   U14708 : OAI222_X1 port map( A1 => n14628, A2 => n16917, B1 => n14564, B2 =>
                           n16914, C1 => n13536, C2 => n16911, ZN => n15321);
   U14709 : OAI222_X1 port map( A1 => n14627, A2 => n16917, B1 => n14563, B2 =>
                           n16914, C1 => n13535, C2 => n16911, ZN => n15304);
   U14710 : OAI222_X1 port map( A1 => n14626, A2 => n16917, B1 => n14562, B2 =>
                           n16914, C1 => n13534, C2 => n16911, ZN => n15287);
   U14711 : OAI222_X1 port map( A1 => n14625, A2 => n16917, B1 => n14561, B2 =>
                           n16914, C1 => n13533, C2 => n16911, ZN => n15270);
   U14712 : OAI222_X1 port map( A1 => n14624, A2 => n16917, B1 => n14560, B2 =>
                           n16914, C1 => n13532, C2 => n16911, ZN => n15253);
   U14713 : OAI222_X1 port map( A1 => n14623, A2 => n16917, B1 => n14559, B2 =>
                           n16914, C1 => n13531, C2 => n16911, ZN => n15236);
   U14714 : OAI222_X1 port map( A1 => n14622, A2 => n16917, B1 => n14558, B2 =>
                           n16914, C1 => n13530, C2 => n16911, ZN => n15187);
   U14715 : OAI222_X1 port map( A1 => n13441, A2 => n16806, B1 => n13377, B2 =>
                           n16803, C1 => n14789, C2 => n16800, ZN => n15917);
   U14716 : OAI222_X1 port map( A1 => n13440, A2 => n16806, B1 => n13376, B2 =>
                           n16803, C1 => n14788, C2 => n16800, ZN => n15900);
   U14717 : OAI222_X1 port map( A1 => n13439, A2 => n16806, B1 => n13375, B2 =>
                           n16803, C1 => n14787, C2 => n16800, ZN => n15883);
   U14718 : OAI222_X1 port map( A1 => n13438, A2 => n16806, B1 => n13374, B2 =>
                           n16803, C1 => n14786, C2 => n16800, ZN => n15866);
   U14719 : OAI222_X1 port map( A1 => n13437, A2 => n16806, B1 => n13373, B2 =>
                           n16803, C1 => n14785, C2 => n16800, ZN => n15849);
   U14720 : OAI222_X1 port map( A1 => n13436, A2 => n16806, B1 => n13372, B2 =>
                           n16803, C1 => n14784, C2 => n16800, ZN => n15832);
   U14721 : OAI222_X1 port map( A1 => n13435, A2 => n16806, B1 => n13371, B2 =>
                           n16803, C1 => n14783, C2 => n16800, ZN => n15815);
   U14722 : OAI222_X1 port map( A1 => n13434, A2 => n16806, B1 => n13370, B2 =>
                           n16803, C1 => n14782, C2 => n16800, ZN => n15766);
   U14723 : OAI222_X1 port map( A1 => n13441, A2 => n16899, B1 => n13377, B2 =>
                           n16896, C1 => n14789, C2 => n16893, ZN => n15336);
   U14724 : OAI222_X1 port map( A1 => n13440, A2 => n16899, B1 => n13376, B2 =>
                           n16896, C1 => n14788, C2 => n16893, ZN => n15319);
   U14725 : OAI222_X1 port map( A1 => n13439, A2 => n16899, B1 => n13375, B2 =>
                           n16896, C1 => n14787, C2 => n16893, ZN => n15302);
   U14726 : OAI222_X1 port map( A1 => n13438, A2 => n16899, B1 => n13374, B2 =>
                           n16896, C1 => n14786, C2 => n16893, ZN => n15285);
   U14727 : OAI222_X1 port map( A1 => n13437, A2 => n16899, B1 => n13373, B2 =>
                           n16896, C1 => n14785, C2 => n16893, ZN => n15268);
   U14728 : OAI222_X1 port map( A1 => n13436, A2 => n16899, B1 => n13372, B2 =>
                           n16896, C1 => n14784, C2 => n16893, ZN => n15251);
   U14729 : OAI222_X1 port map( A1 => n13435, A2 => n16899, B1 => n13371, B2 =>
                           n16896, C1 => n14783, C2 => n16893, ZN => n15234);
   U14730 : OAI222_X1 port map( A1 => n13434, A2 => n16899, B1 => n13370, B2 =>
                           n16896, C1 => n14782, C2 => n16893, ZN => n15185);
   U14731 : OAI222_X1 port map( A1 => n13465, A2 => n16804, B1 => n13401, B2 =>
                           n16801, C1 => n14813, C2 => n16798, ZN => n16325);
   U14732 : OAI222_X1 port map( A1 => n13464, A2 => n16804, B1 => n13400, B2 =>
                           n16801, C1 => n14812, C2 => n16798, ZN => n16308);
   U14733 : OAI222_X1 port map( A1 => n13463, A2 => n16804, B1 => n13399, B2 =>
                           n16801, C1 => n14811, C2 => n16798, ZN => n16291);
   U14734 : OAI222_X1 port map( A1 => n13462, A2 => n16804, B1 => n13398, B2 =>
                           n16801, C1 => n14810, C2 => n16798, ZN => n16274);
   U14735 : OAI222_X1 port map( A1 => n13461, A2 => n16804, B1 => n13397, B2 =>
                           n16801, C1 => n14809, C2 => n16798, ZN => n16257);
   U14736 : OAI222_X1 port map( A1 => n13460, A2 => n16804, B1 => n13396, B2 =>
                           n16801, C1 => n14808, C2 => n16798, ZN => n16240);
   U14737 : OAI222_X1 port map( A1 => n13459, A2 => n16804, B1 => n13395, B2 =>
                           n16801, C1 => n14807, C2 => n16798, ZN => n16223);
   U14738 : OAI222_X1 port map( A1 => n13458, A2 => n16804, B1 => n13394, B2 =>
                           n16801, C1 => n14806, C2 => n16798, ZN => n16206);
   U14739 : OAI222_X1 port map( A1 => n13457, A2 => n16804, B1 => n13393, B2 =>
                           n16801, C1 => n14805, C2 => n16798, ZN => n16189);
   U14740 : OAI222_X1 port map( A1 => n13456, A2 => n16804, B1 => n13392, B2 =>
                           n16801, C1 => n14804, C2 => n16798, ZN => n16172);
   U14741 : OAI222_X1 port map( A1 => n13455, A2 => n16804, B1 => n13391, B2 =>
                           n16801, C1 => n14803, C2 => n16798, ZN => n16155);
   U14742 : OAI222_X1 port map( A1 => n13454, A2 => n16804, B1 => n13390, B2 =>
                           n16801, C1 => n14802, C2 => n16798, ZN => n16138);
   U14743 : OAI222_X1 port map( A1 => n13453, A2 => n16805, B1 => n13389, B2 =>
                           n16802, C1 => n14801, C2 => n16799, ZN => n16121);
   U14744 : OAI222_X1 port map( A1 => n13452, A2 => n16805, B1 => n13388, B2 =>
                           n16802, C1 => n14800, C2 => n16799, ZN => n16104);
   U14745 : OAI222_X1 port map( A1 => n13451, A2 => n16805, B1 => n13387, B2 =>
                           n16802, C1 => n14799, C2 => n16799, ZN => n16087);
   U14746 : OAI222_X1 port map( A1 => n13450, A2 => n16805, B1 => n13386, B2 =>
                           n16802, C1 => n14798, C2 => n16799, ZN => n16070);
   U14747 : OAI222_X1 port map( A1 => n13449, A2 => n16805, B1 => n13385, B2 =>
                           n16802, C1 => n14797, C2 => n16799, ZN => n16053);
   U14748 : OAI222_X1 port map( A1 => n13448, A2 => n16805, B1 => n13384, B2 =>
                           n16802, C1 => n14796, C2 => n16799, ZN => n16036);
   U14749 : OAI222_X1 port map( A1 => n13447, A2 => n16805, B1 => n13383, B2 =>
                           n16802, C1 => n14795, C2 => n16799, ZN => n16019);
   U14750 : OAI222_X1 port map( A1 => n13446, A2 => n16805, B1 => n13382, B2 =>
                           n16802, C1 => n14794, C2 => n16799, ZN => n16002);
   U14751 : OAI222_X1 port map( A1 => n13445, A2 => n16805, B1 => n13381, B2 =>
                           n16802, C1 => n14793, C2 => n16799, ZN => n15985);
   U14752 : OAI222_X1 port map( A1 => n13444, A2 => n16805, B1 => n13380, B2 =>
                           n16802, C1 => n14792, C2 => n16799, ZN => n15968);
   U14753 : OAI222_X1 port map( A1 => n13443, A2 => n16805, B1 => n13379, B2 =>
                           n16802, C1 => n14791, C2 => n16799, ZN => n15951);
   U14754 : OAI222_X1 port map( A1 => n13442, A2 => n16805, B1 => n13378, B2 =>
                           n16802, C1 => n14790, C2 => n16799, ZN => n15934);
   U14755 : OAI222_X1 port map( A1 => n13465, A2 => n16897, B1 => n13401, B2 =>
                           n16894, C1 => n14813, C2 => n16891, ZN => n15744);
   U14756 : OAI222_X1 port map( A1 => n13464, A2 => n16897, B1 => n13400, B2 =>
                           n16894, C1 => n14812, C2 => n16891, ZN => n15727);
   U14757 : OAI222_X1 port map( A1 => n13463, A2 => n16897, B1 => n13399, B2 =>
                           n16894, C1 => n14811, C2 => n16891, ZN => n15710);
   U14758 : OAI222_X1 port map( A1 => n13462, A2 => n16897, B1 => n13398, B2 =>
                           n16894, C1 => n14810, C2 => n16891, ZN => n15693);
   U14759 : OAI222_X1 port map( A1 => n13461, A2 => n16897, B1 => n13397, B2 =>
                           n16894, C1 => n14809, C2 => n16891, ZN => n15676);
   U14760 : OAI222_X1 port map( A1 => n13460, A2 => n16897, B1 => n13396, B2 =>
                           n16894, C1 => n14808, C2 => n16891, ZN => n15659);
   U14761 : OAI222_X1 port map( A1 => n13459, A2 => n16897, B1 => n13395, B2 =>
                           n16894, C1 => n14807, C2 => n16891, ZN => n15642);
   U14762 : OAI222_X1 port map( A1 => n13458, A2 => n16897, B1 => n13394, B2 =>
                           n16894, C1 => n14806, C2 => n16891, ZN => n15625);
   U14763 : OAI222_X1 port map( A1 => n13457, A2 => n16897, B1 => n13393, B2 =>
                           n16894, C1 => n14805, C2 => n16891, ZN => n15608);
   U14764 : OAI222_X1 port map( A1 => n13456, A2 => n16897, B1 => n13392, B2 =>
                           n16894, C1 => n14804, C2 => n16891, ZN => n15591);
   U14765 : OAI222_X1 port map( A1 => n13455, A2 => n16897, B1 => n13391, B2 =>
                           n16894, C1 => n14803, C2 => n16891, ZN => n15574);
   U14766 : OAI222_X1 port map( A1 => n13454, A2 => n16897, B1 => n13390, B2 =>
                           n16894, C1 => n14802, C2 => n16891, ZN => n15557);
   U14767 : OAI222_X1 port map( A1 => n13453, A2 => n16898, B1 => n13389, B2 =>
                           n16895, C1 => n14801, C2 => n16892, ZN => n15540);
   U14768 : OAI222_X1 port map( A1 => n13452, A2 => n16898, B1 => n13388, B2 =>
                           n16895, C1 => n14800, C2 => n16892, ZN => n15523);
   U14769 : OAI222_X1 port map( A1 => n13451, A2 => n16898, B1 => n13387, B2 =>
                           n16895, C1 => n14799, C2 => n16892, ZN => n15506);
   U14770 : OAI222_X1 port map( A1 => n13450, A2 => n16898, B1 => n13386, B2 =>
                           n16895, C1 => n14798, C2 => n16892, ZN => n15489);
   U14771 : OAI222_X1 port map( A1 => n13449, A2 => n16898, B1 => n13385, B2 =>
                           n16895, C1 => n14797, C2 => n16892, ZN => n15472);
   U14772 : OAI222_X1 port map( A1 => n13448, A2 => n16898, B1 => n13384, B2 =>
                           n16895, C1 => n14796, C2 => n16892, ZN => n15455);
   U14773 : OAI222_X1 port map( A1 => n13447, A2 => n16898, B1 => n13383, B2 =>
                           n16895, C1 => n14795, C2 => n16892, ZN => n15438);
   U14774 : OAI222_X1 port map( A1 => n13446, A2 => n16898, B1 => n13382, B2 =>
                           n16895, C1 => n14794, C2 => n16892, ZN => n15421);
   U14775 : OAI222_X1 port map( A1 => n13445, A2 => n16898, B1 => n13381, B2 =>
                           n16895, C1 => n14793, C2 => n16892, ZN => n15404);
   U14776 : OAI222_X1 port map( A1 => n13444, A2 => n16898, B1 => n13380, B2 =>
                           n16895, C1 => n14792, C2 => n16892, ZN => n15387);
   U14777 : OAI222_X1 port map( A1 => n13443, A2 => n16898, B1 => n13379, B2 =>
                           n16895, C1 => n14791, C2 => n16892, ZN => n15370);
   U14778 : OAI222_X1 port map( A1 => n13442, A2 => n16898, B1 => n13378, B2 =>
                           n16895, C1 => n14790, C2 => n16892, ZN => n15353);
   U14779 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_0_port, C1 => n16751, 
                           C2 => n16510, A => n16337, ZN => n16320);
   U14780 : AOI21_X1 port map( B1 => n16338, B2 => n16339, A => n16748, ZN => 
                           n16337);
   U14781 : AOI221_X1 port map( B1 => n16735, B2 => n15052, C1 => n16734, C2 =>
                           n15100, A => n16341, ZN => n16338);
   U14782 : AOI221_X1 port map( B1 => n16745, B2 => n15028, C1 => n16742, C2 =>
                           n15076, A => n16340, ZN => n16339);
   U14783 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_1_port, C1 => n16751, 
                           C2 => n16511, A => n16315, ZN => n16303);
   U14784 : AOI21_X1 port map( B1 => n16316, B2 => n16317, A => n16748, ZN => 
                           n16315);
   U14785 : AOI221_X1 port map( B1 => n16737, B2 => n15051, C1 => n16734, C2 =>
                           n15099, A => n16319, ZN => n16316);
   U14786 : AOI221_X1 port map( B1 => n16747, B2 => n15027, C1 => n16744, C2 =>
                           n15075, A => n16318, ZN => n16317);
   U14787 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_2_port, C1 => n16751, 
                           C2 => n16512, A => n16298, ZN => n16286);
   U14788 : AOI21_X1 port map( B1 => n16299, B2 => n16300, A => n16748, ZN => 
                           n16298);
   U14789 : AOI221_X1 port map( B1 => n16737, B2 => n15050, C1 => n16734, C2 =>
                           n15098, A => n16302, ZN => n16299);
   U14790 : AOI221_X1 port map( B1 => n16747, B2 => n15026, C1 => n16744, C2 =>
                           n15074, A => n16301, ZN => n16300);
   U14791 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_3_port, C1 => n16751, 
                           C2 => n16513, A => n16281, ZN => n16269);
   U14792 : AOI21_X1 port map( B1 => n16282, B2 => n16283, A => n16748, ZN => 
                           n16281);
   U14793 : AOI221_X1 port map( B1 => n16737, B2 => n15049, C1 => n16734, C2 =>
                           n15097, A => n16285, ZN => n16282);
   U14794 : AOI221_X1 port map( B1 => n16747, B2 => n15025, C1 => n16744, C2 =>
                           n15073, A => n16284, ZN => n16283);
   U14795 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_4_port, C1 => n16751, 
                           C2 => n16514, A => n16264, ZN => n16252);
   U14796 : AOI21_X1 port map( B1 => n16265, B2 => n16266, A => n16748, ZN => 
                           n16264);
   U14797 : AOI221_X1 port map( B1 => n16737, B2 => n15048, C1 => n16734, C2 =>
                           n15096, A => n16268, ZN => n16265);
   U14798 : AOI221_X1 port map( B1 => n16747, B2 => n15024, C1 => n16744, C2 =>
                           n15072, A => n16267, ZN => n16266);
   U14799 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_5_port, C1 => n16751, 
                           C2 => n16515, A => n16247, ZN => n16235);
   U14800 : AOI21_X1 port map( B1 => n16248, B2 => n16249, A => n16748, ZN => 
                           n16247);
   U14801 : AOI221_X1 port map( B1 => n16737, B2 => n15047, C1 => n16734, C2 =>
                           n15095, A => n16251, ZN => n16248);
   U14802 : AOI221_X1 port map( B1 => n16747, B2 => n15023, C1 => n16744, C2 =>
                           n15071, A => n16250, ZN => n16249);
   U14803 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_6_port, C1 => n16751, 
                           C2 => n16516, A => n16230, ZN => n16218);
   U14804 : AOI21_X1 port map( B1 => n16231, B2 => n16232, A => n16748, ZN => 
                           n16230);
   U14805 : AOI221_X1 port map( B1 => n16737, B2 => n15046, C1 => n16734, C2 =>
                           n15094, A => n16234, ZN => n16231);
   U14806 : AOI221_X1 port map( B1 => n16747, B2 => n15022, C1 => n16744, C2 =>
                           n15070, A => n16233, ZN => n16232);
   U14807 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_7_port, C1 => n16751, 
                           C2 => n16517, A => n16213, ZN => n16201);
   U14808 : AOI21_X1 port map( B1 => n16214, B2 => n16215, A => n16748, ZN => 
                           n16213);
   U14809 : AOI221_X1 port map( B1 => n16737, B2 => n15045, C1 => n16734, C2 =>
                           n15093, A => n16217, ZN => n16214);
   U14810 : AOI221_X1 port map( B1 => n16747, B2 => n15021, C1 => n16744, C2 =>
                           n15069, A => n16216, ZN => n16215);
   U14811 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_8_port, C1 => n16751, 
                           C2 => n16518, A => n16196, ZN => n16184);
   U14812 : AOI21_X1 port map( B1 => n16197, B2 => n16198, A => n16748, ZN => 
                           n16196);
   U14813 : AOI221_X1 port map( B1 => n16737, B2 => n15044, C1 => n16733, C2 =>
                           n15092, A => n16200, ZN => n16197);
   U14814 : AOI221_X1 port map( B1 => n16747, B2 => n15020, C1 => n16744, C2 =>
                           n15068, A => n16199, ZN => n16198);
   U14815 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_9_port, C1 => n16751, 
                           C2 => n16519, A => n16179, ZN => n16167);
   U14816 : AOI21_X1 port map( B1 => n16180, B2 => n16181, A => n16748, ZN => 
                           n16179);
   U14817 : AOI221_X1 port map( B1 => n16736, B2 => n15043, C1 => n16733, C2 =>
                           n15091, A => n16183, ZN => n16180);
   U14818 : AOI221_X1 port map( B1 => n16746, B2 => n15019, C1 => n16743, C2 =>
                           n15067, A => n16182, ZN => n16181);
   U14819 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_10_port, C1 => n16751,
                           C2 => n16520, A => n16162, ZN => n16150);
   U14820 : AOI21_X1 port map( B1 => n16163, B2 => n16164, A => n16748, ZN => 
                           n16162);
   U14821 : AOI221_X1 port map( B1 => n16736, B2 => n15042, C1 => n16733, C2 =>
                           n15090, A => n16166, ZN => n16163);
   U14822 : AOI221_X1 port map( B1 => n16746, B2 => n15018, C1 => n16743, C2 =>
                           n15066, A => n16165, ZN => n16164);
   U14823 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_11_port, C1 => n16751,
                           C2 => n16521, A => n16145, ZN => n16133);
   U14824 : AOI21_X1 port map( B1 => n16146, B2 => n16147, A => n16748, ZN => 
                           n16145);
   U14825 : AOI221_X1 port map( B1 => n16736, B2 => n15041, C1 => n16733, C2 =>
                           n15089, A => n16149, ZN => n16146);
   U14826 : AOI221_X1 port map( B1 => n16746, B2 => n15017, C1 => n16743, C2 =>
                           n15065, A => n16148, ZN => n16147);
   U14827 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_12_port, C1 => n16752,
                           C2 => n16522, A => n16128, ZN => n16116);
   U14828 : AOI21_X1 port map( B1 => n16129, B2 => n16130, A => n16749, ZN => 
                           n16128);
   U14829 : AOI221_X1 port map( B1 => n16736, B2 => n15040, C1 => n16733, C2 =>
                           n15088, A => n16132, ZN => n16129);
   U14830 : AOI221_X1 port map( B1 => n16746, B2 => n15016, C1 => n16743, C2 =>
                           n15064, A => n16131, ZN => n16130);
   U14831 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_13_port, C1 => n16752,
                           C2 => n16523, A => n16111, ZN => n16099);
   U14832 : AOI21_X1 port map( B1 => n16112, B2 => n16113, A => n16749, ZN => 
                           n16111);
   U14833 : AOI221_X1 port map( B1 => n16736, B2 => n15039, C1 => n16733, C2 =>
                           n15087, A => n16115, ZN => n16112);
   U14834 : AOI221_X1 port map( B1 => n16746, B2 => n15015, C1 => n16743, C2 =>
                           n15063, A => n16114, ZN => n16113);
   U14835 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_14_port, C1 => n16752,
                           C2 => n16524, A => n16094, ZN => n16082);
   U14836 : AOI21_X1 port map( B1 => n16095, B2 => n16096, A => n16749, ZN => 
                           n16094);
   U14837 : AOI221_X1 port map( B1 => n16736, B2 => n15038, C1 => n16733, C2 =>
                           n15086, A => n16098, ZN => n16095);
   U14838 : AOI221_X1 port map( B1 => n16746, B2 => n15014, C1 => n16743, C2 =>
                           n15062, A => n16097, ZN => n16096);
   U14839 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_15_port, C1 => n16752,
                           C2 => n16525, A => n16077, ZN => n16065);
   U14840 : AOI21_X1 port map( B1 => n16078, B2 => n16079, A => n16749, ZN => 
                           n16077);
   U14841 : AOI221_X1 port map( B1 => n16736, B2 => n15037, C1 => n16733, C2 =>
                           n15085, A => n16081, ZN => n16078);
   U14842 : AOI221_X1 port map( B1 => n16746, B2 => n15013, C1 => n16743, C2 =>
                           n15061, A => n16080, ZN => n16079);
   U14843 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_16_port, C1 => n16752,
                           C2 => n16526, A => n16060, ZN => n16048);
   U14844 : AOI21_X1 port map( B1 => n16061, B2 => n16062, A => n16749, ZN => 
                           n16060);
   U14845 : AOI221_X1 port map( B1 => n16736, B2 => n15036, C1 => n16733, C2 =>
                           n15084, A => n16064, ZN => n16061);
   U14846 : AOI221_X1 port map( B1 => n16746, B2 => n15012, C1 => n16743, C2 =>
                           n15060, A => n16063, ZN => n16062);
   U14847 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_17_port, C1 => n16752,
                           C2 => n16527, A => n16043, ZN => n16031);
   U14848 : AOI21_X1 port map( B1 => n16044, B2 => n16045, A => n16749, ZN => 
                           n16043);
   U14849 : AOI221_X1 port map( B1 => n16736, B2 => n15035, C1 => n16733, C2 =>
                           n15083, A => n16047, ZN => n16044);
   U14850 : AOI221_X1 port map( B1 => n16746, B2 => n15011, C1 => n16743, C2 =>
                           n15059, A => n16046, ZN => n16045);
   U14851 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_18_port, C1 => n16752,
                           C2 => n16528, A => n16026, ZN => n16014);
   U14852 : AOI21_X1 port map( B1 => n16027, B2 => n16028, A => n16749, ZN => 
                           n16026);
   U14853 : AOI221_X1 port map( B1 => n16736, B2 => n15034, C1 => n16733, C2 =>
                           n15082, A => n16030, ZN => n16027);
   U14854 : AOI221_X1 port map( B1 => n16746, B2 => n15010, C1 => n16743, C2 =>
                           n15058, A => n16029, ZN => n16028);
   U14855 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_19_port, C1 => n16752,
                           C2 => n16529, A => n16009, ZN => n15997);
   U14856 : AOI21_X1 port map( B1 => n16010, B2 => n16011, A => n16749, ZN => 
                           n16009);
   U14857 : AOI221_X1 port map( B1 => n16736, B2 => n15033, C1 => n16732, C2 =>
                           n15081, A => n16013, ZN => n16010);
   U14858 : AOI221_X1 port map( B1 => n16746, B2 => n15009, C1 => n16743, C2 =>
                           n15057, A => n16012, ZN => n16011);
   U14859 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_20_port, C1 => n16752,
                           C2 => n16530, A => n15992, ZN => n15980);
   U14860 : AOI21_X1 port map( B1 => n15993, B2 => n15994, A => n16749, ZN => 
                           n15992);
   U14861 : AOI221_X1 port map( B1 => n16735, B2 => n15032, C1 => n16732, C2 =>
                           n15080, A => n15996, ZN => n15993);
   U14862 : AOI221_X1 port map( B1 => n16745, B2 => n15008, C1 => n16742, C2 =>
                           n15056, A => n15995, ZN => n15994);
   U14863 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_21_port, C1 => n16752,
                           C2 => n16531, A => n15975, ZN => n15963);
   U14864 : AOI21_X1 port map( B1 => n15976, B2 => n15977, A => n16749, ZN => 
                           n15975);
   U14865 : AOI221_X1 port map( B1 => n16735, B2 => n15031, C1 => n16732, C2 =>
                           n15079, A => n15979, ZN => n15976);
   U14866 : AOI221_X1 port map( B1 => n16745, B2 => n15007, C1 => n16742, C2 =>
                           n15055, A => n15978, ZN => n15977);
   U14867 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_22_port, C1 => n16752,
                           C2 => n16532, A => n15958, ZN => n15946);
   U14868 : AOI21_X1 port map( B1 => n15959, B2 => n15960, A => n16749, ZN => 
                           n15958);
   U14869 : AOI221_X1 port map( B1 => n16735, B2 => n15030, C1 => n16732, C2 =>
                           n15078, A => n15962, ZN => n15959);
   U14870 : AOI221_X1 port map( B1 => n16745, B2 => n15006, C1 => n16742, C2 =>
                           n15054, A => n15961, ZN => n15960);
   U14871 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_23_port, C1 => n16752,
                           C2 => n16533, A => n15941, ZN => n15929);
   U14872 : AOI21_X1 port map( B1 => n15942, B2 => n15943, A => n16749, ZN => 
                           n15941);
   U14873 : AOI221_X1 port map( B1 => n16735, B2 => n15029, C1 => n16732, C2 =>
                           n15077, A => n15945, ZN => n15942);
   U14874 : AOI221_X1 port map( B1 => n16745, B2 => n15005, C1 => n16742, C2 =>
                           n15053, A => n15944, ZN => n15943);
   U14875 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_0_port, C1 => n16844, 
                           C2 => n16510, A => n15756, ZN => n15739);
   U14876 : AOI21_X1 port map( B1 => n15757, B2 => n15758, A => n16841, ZN => 
                           n15756);
   U14877 : AOI221_X1 port map( B1 => n16828, B2 => n15052, C1 => n16827, C2 =>
                           n15100, A => n15760, ZN => n15757);
   U14878 : AOI221_X1 port map( B1 => n16838, B2 => n15028, C1 => n16835, C2 =>
                           n15076, A => n15759, ZN => n15758);
   U14879 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_1_port, C1 => n16844, 
                           C2 => n16511, A => n15734, ZN => n15722);
   U14880 : AOI21_X1 port map( B1 => n15735, B2 => n15736, A => n16841, ZN => 
                           n15734);
   U14881 : AOI221_X1 port map( B1 => n16830, B2 => n15051, C1 => n16827, C2 =>
                           n15099, A => n15738, ZN => n15735);
   U14882 : AOI221_X1 port map( B1 => n16840, B2 => n15027, C1 => n16837, C2 =>
                           n15075, A => n15737, ZN => n15736);
   U14883 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_2_port, C1 => n16844, 
                           C2 => n16512, A => n15717, ZN => n15705);
   U14884 : AOI21_X1 port map( B1 => n15718, B2 => n15719, A => n16841, ZN => 
                           n15717);
   U14885 : AOI221_X1 port map( B1 => n16830, B2 => n15050, C1 => n16827, C2 =>
                           n15098, A => n15721, ZN => n15718);
   U14886 : AOI221_X1 port map( B1 => n16840, B2 => n15026, C1 => n16837, C2 =>
                           n15074, A => n15720, ZN => n15719);
   U14887 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_3_port, C1 => n16844, 
                           C2 => n16513, A => n15700, ZN => n15688);
   U14888 : AOI21_X1 port map( B1 => n15701, B2 => n15702, A => n16841, ZN => 
                           n15700);
   U14889 : AOI221_X1 port map( B1 => n16830, B2 => n15049, C1 => n16827, C2 =>
                           n15097, A => n15704, ZN => n15701);
   U14890 : AOI221_X1 port map( B1 => n16840, B2 => n15025, C1 => n16837, C2 =>
                           n15073, A => n15703, ZN => n15702);
   U14891 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_4_port, C1 => n16844, 
                           C2 => n16514, A => n15683, ZN => n15671);
   U14892 : AOI21_X1 port map( B1 => n15684, B2 => n15685, A => n16841, ZN => 
                           n15683);
   U14893 : AOI221_X1 port map( B1 => n16830, B2 => n15048, C1 => n16827, C2 =>
                           n15096, A => n15687, ZN => n15684);
   U14894 : AOI221_X1 port map( B1 => n16840, B2 => n15024, C1 => n16837, C2 =>
                           n15072, A => n15686, ZN => n15685);
   U14895 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_5_port, C1 => n16844, 
                           C2 => n16515, A => n15666, ZN => n15654);
   U14896 : AOI21_X1 port map( B1 => n15667, B2 => n15668, A => n16841, ZN => 
                           n15666);
   U14897 : AOI221_X1 port map( B1 => n16830, B2 => n15047, C1 => n16827, C2 =>
                           n15095, A => n15670, ZN => n15667);
   U14898 : AOI221_X1 port map( B1 => n16840, B2 => n15023, C1 => n16837, C2 =>
                           n15071, A => n15669, ZN => n15668);
   U14899 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_6_port, C1 => n16844, 
                           C2 => n16516, A => n15649, ZN => n15637);
   U14900 : AOI21_X1 port map( B1 => n15650, B2 => n15651, A => n16841, ZN => 
                           n15649);
   U14901 : AOI221_X1 port map( B1 => n16830, B2 => n15046, C1 => n16827, C2 =>
                           n15094, A => n15653, ZN => n15650);
   U14902 : AOI221_X1 port map( B1 => n16840, B2 => n15022, C1 => n16837, C2 =>
                           n15070, A => n15652, ZN => n15651);
   U14903 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_7_port, C1 => n16844, 
                           C2 => n16517, A => n15632, ZN => n15620);
   U14904 : AOI21_X1 port map( B1 => n15633, B2 => n15634, A => n16841, ZN => 
                           n15632);
   U14905 : AOI221_X1 port map( B1 => n16830, B2 => n15045, C1 => n16827, C2 =>
                           n15093, A => n15636, ZN => n15633);
   U14906 : AOI221_X1 port map( B1 => n16840, B2 => n15021, C1 => n16837, C2 =>
                           n15069, A => n15635, ZN => n15634);
   U14907 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_8_port, C1 => n16844, 
                           C2 => n16518, A => n15615, ZN => n15603);
   U14908 : AOI21_X1 port map( B1 => n15616, B2 => n15617, A => n16841, ZN => 
                           n15615);
   U14909 : AOI221_X1 port map( B1 => n16830, B2 => n15044, C1 => n16826, C2 =>
                           n15092, A => n15619, ZN => n15616);
   U14910 : AOI221_X1 port map( B1 => n16840, B2 => n15020, C1 => n16837, C2 =>
                           n15068, A => n15618, ZN => n15617);
   U14911 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_9_port, C1 => n16844, 
                           C2 => n16519, A => n15598, ZN => n15586);
   U14912 : AOI21_X1 port map( B1 => n15599, B2 => n15600, A => n16841, ZN => 
                           n15598);
   U14913 : AOI221_X1 port map( B1 => n16829, B2 => n15043, C1 => n16826, C2 =>
                           n15091, A => n15602, ZN => n15599);
   U14914 : AOI221_X1 port map( B1 => n16839, B2 => n15019, C1 => n16836, C2 =>
                           n15067, A => n15601, ZN => n15600);
   U14915 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_10_port, C1 => n16844,
                           C2 => n16520, A => n15581, ZN => n15569);
   U14916 : AOI21_X1 port map( B1 => n15582, B2 => n15583, A => n16841, ZN => 
                           n15581);
   U14917 : AOI221_X1 port map( B1 => n16829, B2 => n15042, C1 => n16826, C2 =>
                           n15090, A => n15585, ZN => n15582);
   U14918 : AOI221_X1 port map( B1 => n16839, B2 => n15018, C1 => n16836, C2 =>
                           n15066, A => n15584, ZN => n15583);
   U14919 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_11_port, C1 => n16844,
                           C2 => n16521, A => n15564, ZN => n15552);
   U14920 : AOI21_X1 port map( B1 => n15565, B2 => n15566, A => n16841, ZN => 
                           n15564);
   U14921 : AOI221_X1 port map( B1 => n16829, B2 => n15041, C1 => n16826, C2 =>
                           n15089, A => n15568, ZN => n15565);
   U14922 : AOI221_X1 port map( B1 => n16839, B2 => n15017, C1 => n16836, C2 =>
                           n15065, A => n15567, ZN => n15566);
   U14923 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_12_port, C1 => n16845,
                           C2 => n16522, A => n15547, ZN => n15535);
   U14924 : AOI21_X1 port map( B1 => n15548, B2 => n15549, A => n16842, ZN => 
                           n15547);
   U14925 : AOI221_X1 port map( B1 => n16829, B2 => n15040, C1 => n16826, C2 =>
                           n15088, A => n15551, ZN => n15548);
   U14926 : AOI221_X1 port map( B1 => n16839, B2 => n15016, C1 => n16836, C2 =>
                           n15064, A => n15550, ZN => n15549);
   U14927 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_13_port, C1 => n16845,
                           C2 => n16523, A => n15530, ZN => n15518);
   U14928 : AOI21_X1 port map( B1 => n15531, B2 => n15532, A => n16842, ZN => 
                           n15530);
   U14929 : AOI221_X1 port map( B1 => n16829, B2 => n15039, C1 => n16826, C2 =>
                           n15087, A => n15534, ZN => n15531);
   U14930 : AOI221_X1 port map( B1 => n16839, B2 => n15015, C1 => n16836, C2 =>
                           n15063, A => n15533, ZN => n15532);
   U14931 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_14_port, C1 => n16845,
                           C2 => n16524, A => n15513, ZN => n15501);
   U14932 : AOI21_X1 port map( B1 => n15514, B2 => n15515, A => n16842, ZN => 
                           n15513);
   U14933 : AOI221_X1 port map( B1 => n16829, B2 => n15038, C1 => n16826, C2 =>
                           n15086, A => n15517, ZN => n15514);
   U14934 : AOI221_X1 port map( B1 => n16839, B2 => n15014, C1 => n16836, C2 =>
                           n15062, A => n15516, ZN => n15515);
   U14935 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_15_port, C1 => n16845,
                           C2 => n16525, A => n15496, ZN => n15484);
   U14936 : AOI21_X1 port map( B1 => n15497, B2 => n15498, A => n16842, ZN => 
                           n15496);
   U14937 : AOI221_X1 port map( B1 => n16829, B2 => n15037, C1 => n16826, C2 =>
                           n15085, A => n15500, ZN => n15497);
   U14938 : AOI221_X1 port map( B1 => n16839, B2 => n15013, C1 => n16836, C2 =>
                           n15061, A => n15499, ZN => n15498);
   U14939 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_16_port, C1 => n16845,
                           C2 => n16526, A => n15479, ZN => n15467);
   U14940 : AOI21_X1 port map( B1 => n15480, B2 => n15481, A => n16842, ZN => 
                           n15479);
   U14941 : AOI221_X1 port map( B1 => n16829, B2 => n15036, C1 => n16826, C2 =>
                           n15084, A => n15483, ZN => n15480);
   U14942 : AOI221_X1 port map( B1 => n16839, B2 => n15012, C1 => n16836, C2 =>
                           n15060, A => n15482, ZN => n15481);
   U14943 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_17_port, C1 => n16845,
                           C2 => n16527, A => n15462, ZN => n15450);
   U14944 : AOI21_X1 port map( B1 => n15463, B2 => n15464, A => n16842, ZN => 
                           n15462);
   U14945 : AOI221_X1 port map( B1 => n16829, B2 => n15035, C1 => n16826, C2 =>
                           n15083, A => n15466, ZN => n15463);
   U14946 : AOI221_X1 port map( B1 => n16839, B2 => n15011, C1 => n16836, C2 =>
                           n15059, A => n15465, ZN => n15464);
   U14947 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_18_port, C1 => n16845,
                           C2 => n16528, A => n15445, ZN => n15433);
   U14948 : AOI21_X1 port map( B1 => n15446, B2 => n15447, A => n16842, ZN => 
                           n15445);
   U14949 : AOI221_X1 port map( B1 => n16829, B2 => n15034, C1 => n16826, C2 =>
                           n15082, A => n15449, ZN => n15446);
   U14950 : AOI221_X1 port map( B1 => n16839, B2 => n15010, C1 => n16836, C2 =>
                           n15058, A => n15448, ZN => n15447);
   U14951 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_19_port, C1 => n16845,
                           C2 => n16529, A => n15428, ZN => n15416);
   U14952 : AOI21_X1 port map( B1 => n15429, B2 => n15430, A => n16842, ZN => 
                           n15428);
   U14953 : AOI221_X1 port map( B1 => n16829, B2 => n15033, C1 => n16825, C2 =>
                           n15081, A => n15432, ZN => n15429);
   U14954 : AOI221_X1 port map( B1 => n16839, B2 => n15009, C1 => n16836, C2 =>
                           n15057, A => n15431, ZN => n15430);
   U14955 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_20_port, C1 => n16845,
                           C2 => n16530, A => n15411, ZN => n15399);
   U14956 : AOI21_X1 port map( B1 => n15412, B2 => n15413, A => n16842, ZN => 
                           n15411);
   U14957 : AOI221_X1 port map( B1 => n16828, B2 => n15032, C1 => n16825, C2 =>
                           n15080, A => n15415, ZN => n15412);
   U14958 : AOI221_X1 port map( B1 => n16838, B2 => n15008, C1 => n16835, C2 =>
                           n15056, A => n15414, ZN => n15413);
   U14959 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_21_port, C1 => n16845,
                           C2 => n16531, A => n15394, ZN => n15382);
   U14960 : AOI21_X1 port map( B1 => n15395, B2 => n15396, A => n16842, ZN => 
                           n15394);
   U14961 : AOI221_X1 port map( B1 => n16828, B2 => n15031, C1 => n16825, C2 =>
                           n15079, A => n15398, ZN => n15395);
   U14962 : AOI221_X1 port map( B1 => n16838, B2 => n15007, C1 => n16835, C2 =>
                           n15055, A => n15397, ZN => n15396);
   U14963 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_22_port, C1 => n16845,
                           C2 => n16532, A => n15377, ZN => n15365);
   U14964 : AOI21_X1 port map( B1 => n15378, B2 => n15379, A => n16842, ZN => 
                           n15377);
   U14965 : AOI221_X1 port map( B1 => n16828, B2 => n15030, C1 => n16825, C2 =>
                           n15078, A => n15381, ZN => n15378);
   U14966 : AOI221_X1 port map( B1 => n16838, B2 => n15006, C1 => n16835, C2 =>
                           n15054, A => n15380, ZN => n15379);
   U14967 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_23_port, C1 => n16845,
                           C2 => n16533, A => n15360, ZN => n15348);
   U14968 : AOI21_X1 port map( B1 => n15361, B2 => n15362, A => n16842, ZN => 
                           n15360);
   U14969 : AOI221_X1 port map( B1 => n16828, B2 => n15029, C1 => n16825, C2 =>
                           n15077, A => n15364, ZN => n15361);
   U14970 : AOI221_X1 port map( B1 => n16838, B2 => n15005, C1 => n16835, C2 =>
                           n15053, A => n15363, ZN => n15362);
   U14971 : OAI221_X1 port map( B1 => n13721, B2 => n16795, C1 => n13433, C2 =>
                           n16792, A => n16332, ZN => n16324);
   U14972 : AOI22_X1 port map( A1 => n16789, A2 => n14932, B1 => n16788, B2 => 
                           n14956, ZN => n16332);
   U14973 : OAI221_X1 port map( B1 => n13720, B2 => n16795, C1 => n13432, C2 =>
                           n16792, A => n16311, ZN => n16307);
   U14974 : AOI22_X1 port map( A1 => n16789, A2 => n14931, B1 => n16788, B2 => 
                           n14955, ZN => n16311);
   U14975 : OAI221_X1 port map( B1 => n13719, B2 => n16795, C1 => n13431, C2 =>
                           n16792, A => n16294, ZN => n16290);
   U14976 : AOI22_X1 port map( A1 => n16789, A2 => n14930, B1 => n16788, B2 => 
                           n14954, ZN => n16294);
   U14977 : OAI221_X1 port map( B1 => n13718, B2 => n16795, C1 => n13430, C2 =>
                           n16792, A => n16277, ZN => n16273);
   U14978 : AOI22_X1 port map( A1 => n16789, A2 => n14929, B1 => n16788, B2 => 
                           n14953, ZN => n16277);
   U14979 : OAI221_X1 port map( B1 => n13717, B2 => n16795, C1 => n13429, C2 =>
                           n16792, A => n16260, ZN => n16256);
   U14980 : AOI22_X1 port map( A1 => n16789, A2 => n14928, B1 => n16788, B2 => 
                           n14952, ZN => n16260);
   U14981 : OAI221_X1 port map( B1 => n13716, B2 => n16795, C1 => n13428, C2 =>
                           n16792, A => n16243, ZN => n16239);
   U14982 : AOI22_X1 port map( A1 => n16789, A2 => n14927, B1 => n16788, B2 => 
                           n14951, ZN => n16243);
   U14983 : OAI221_X1 port map( B1 => n13715, B2 => n16795, C1 => n13427, C2 =>
                           n16792, A => n16226, ZN => n16222);
   U14984 : AOI22_X1 port map( A1 => n16789, A2 => n14926, B1 => n16788, B2 => 
                           n14950, ZN => n16226);
   U14985 : OAI221_X1 port map( B1 => n13714, B2 => n16795, C1 => n13426, C2 =>
                           n16792, A => n16209, ZN => n16205);
   U14986 : AOI22_X1 port map( A1 => n16789, A2 => n14925, B1 => n16788, B2 => 
                           n14949, ZN => n16209);
   U14987 : OAI221_X1 port map( B1 => n13713, B2 => n16795, C1 => n13425, C2 =>
                           n16792, A => n16192, ZN => n16188);
   U14988 : AOI22_X1 port map( A1 => n16789, A2 => n14924, B1 => n16787, B2 => 
                           n14948, ZN => n16192);
   U14989 : OAI221_X1 port map( B1 => n13712, B2 => n16795, C1 => n13424, C2 =>
                           n16792, A => n16175, ZN => n16171);
   U14990 : AOI22_X1 port map( A1 => n16789, A2 => n14923, B1 => n16787, B2 => 
                           n14947, ZN => n16175);
   U14991 : OAI221_X1 port map( B1 => n13711, B2 => n16795, C1 => n13423, C2 =>
                           n16792, A => n16158, ZN => n16154);
   U14992 : AOI22_X1 port map( A1 => n16789, A2 => n14922, B1 => n16787, B2 => 
                           n14946, ZN => n16158);
   U14993 : OAI221_X1 port map( B1 => n13710, B2 => n16795, C1 => n13422, C2 =>
                           n16792, A => n16141, ZN => n16137);
   U14994 : AOI22_X1 port map( A1 => n16789, A2 => n14921, B1 => n16787, B2 => 
                           n14945, ZN => n16141);
   U14995 : OAI221_X1 port map( B1 => n13709, B2 => n16796, C1 => n13421, C2 =>
                           n16793, A => n16124, ZN => n16120);
   U14996 : AOI22_X1 port map( A1 => n16790, A2 => n14920, B1 => n16787, B2 => 
                           n14944, ZN => n16124);
   U14997 : OAI221_X1 port map( B1 => n13708, B2 => n16796, C1 => n13420, C2 =>
                           n16793, A => n16107, ZN => n16103);
   U14998 : AOI22_X1 port map( A1 => n16790, A2 => n14919, B1 => n16787, B2 => 
                           n14943, ZN => n16107);
   U14999 : OAI221_X1 port map( B1 => n13707, B2 => n16796, C1 => n13419, C2 =>
                           n16793, A => n16090, ZN => n16086);
   U15000 : AOI22_X1 port map( A1 => n16790, A2 => n14918, B1 => n16787, B2 => 
                           n14942, ZN => n16090);
   U15001 : OAI221_X1 port map( B1 => n13706, B2 => n16796, C1 => n13418, C2 =>
                           n16793, A => n16073, ZN => n16069);
   U15002 : AOI22_X1 port map( A1 => n16790, A2 => n14917, B1 => n16787, B2 => 
                           n14941, ZN => n16073);
   U15003 : OAI221_X1 port map( B1 => n13705, B2 => n16796, C1 => n13417, C2 =>
                           n16793, A => n16056, ZN => n16052);
   U15004 : AOI22_X1 port map( A1 => n16790, A2 => n14916, B1 => n16787, B2 => 
                           n14940, ZN => n16056);
   U15005 : OAI221_X1 port map( B1 => n13704, B2 => n16796, C1 => n13416, C2 =>
                           n16793, A => n16039, ZN => n16035);
   U15006 : AOI22_X1 port map( A1 => n16790, A2 => n14915, B1 => n16787, B2 => 
                           n14939, ZN => n16039);
   U15007 : OAI221_X1 port map( B1 => n13703, B2 => n16796, C1 => n13415, C2 =>
                           n16793, A => n16022, ZN => n16018);
   U15008 : AOI22_X1 port map( A1 => n16790, A2 => n14914, B1 => n16787, B2 => 
                           n14938, ZN => n16022);
   U15009 : OAI221_X1 port map( B1 => n13702, B2 => n16796, C1 => n13414, C2 =>
                           n16793, A => n16005, ZN => n16001);
   U15010 : AOI22_X1 port map( A1 => n16790, A2 => n14913, B1 => n16787, B2 => 
                           n14937, ZN => n16005);
   U15011 : OAI221_X1 port map( B1 => n13701, B2 => n16796, C1 => n13413, C2 =>
                           n16793, A => n15988, ZN => n15984);
   U15012 : AOI22_X1 port map( A1 => n16790, A2 => n14912, B1 => n16786, B2 => 
                           n14936, ZN => n15988);
   U15013 : OAI221_X1 port map( B1 => n13700, B2 => n16796, C1 => n13412, C2 =>
                           n16793, A => n15971, ZN => n15967);
   U15014 : AOI22_X1 port map( A1 => n16790, A2 => n14911, B1 => n16786, B2 => 
                           n14935, ZN => n15971);
   U15015 : OAI221_X1 port map( B1 => n13699, B2 => n16796, C1 => n13411, C2 =>
                           n16793, A => n15954, ZN => n15950);
   U15016 : AOI22_X1 port map( A1 => n16790, A2 => n14910, B1 => n16786, B2 => 
                           n14934, ZN => n15954);
   U15017 : OAI221_X1 port map( B1 => n13698, B2 => n16796, C1 => n13410, C2 =>
                           n16793, A => n15937, ZN => n15933);
   U15018 : AOI22_X1 port map( A1 => n16790, A2 => n14909, B1 => n16786, B2 => 
                           n14933, ZN => n15937);
   U15019 : OAI221_X1 port map( B1 => n13721, B2 => n16888, C1 => n13433, C2 =>
                           n16885, A => n15751, ZN => n15743);
   U15020 : AOI22_X1 port map( A1 => n16882, A2 => n14932, B1 => n16881, B2 => 
                           n14956, ZN => n15751);
   U15021 : OAI221_X1 port map( B1 => n13720, B2 => n16888, C1 => n13432, C2 =>
                           n16885, A => n15730, ZN => n15726);
   U15022 : AOI22_X1 port map( A1 => n16882, A2 => n14931, B1 => n16881, B2 => 
                           n14955, ZN => n15730);
   U15023 : OAI221_X1 port map( B1 => n13719, B2 => n16888, C1 => n13431, C2 =>
                           n16885, A => n15713, ZN => n15709);
   U15024 : AOI22_X1 port map( A1 => n16882, A2 => n14930, B1 => n16881, B2 => 
                           n14954, ZN => n15713);
   U15025 : OAI221_X1 port map( B1 => n13718, B2 => n16888, C1 => n13430, C2 =>
                           n16885, A => n15696, ZN => n15692);
   U15026 : AOI22_X1 port map( A1 => n16882, A2 => n14929, B1 => n16881, B2 => 
                           n14953, ZN => n15696);
   U15027 : OAI221_X1 port map( B1 => n13717, B2 => n16888, C1 => n13429, C2 =>
                           n16885, A => n15679, ZN => n15675);
   U15028 : AOI22_X1 port map( A1 => n16882, A2 => n14928, B1 => n16881, B2 => 
                           n14952, ZN => n15679);
   U15029 : OAI221_X1 port map( B1 => n13716, B2 => n16888, C1 => n13428, C2 =>
                           n16885, A => n15662, ZN => n15658);
   U15030 : AOI22_X1 port map( A1 => n16882, A2 => n14927, B1 => n16881, B2 => 
                           n14951, ZN => n15662);
   U15031 : OAI221_X1 port map( B1 => n13715, B2 => n16888, C1 => n13427, C2 =>
                           n16885, A => n15645, ZN => n15641);
   U15032 : AOI22_X1 port map( A1 => n16882, A2 => n14926, B1 => n16881, B2 => 
                           n14950, ZN => n15645);
   U15033 : OAI221_X1 port map( B1 => n13714, B2 => n16888, C1 => n13426, C2 =>
                           n16885, A => n15628, ZN => n15624);
   U15034 : AOI22_X1 port map( A1 => n16882, A2 => n14925, B1 => n16881, B2 => 
                           n14949, ZN => n15628);
   U15035 : OAI221_X1 port map( B1 => n13713, B2 => n16888, C1 => n13425, C2 =>
                           n16885, A => n15611, ZN => n15607);
   U15036 : AOI22_X1 port map( A1 => n16882, A2 => n14924, B1 => n16880, B2 => 
                           n14948, ZN => n15611);
   U15037 : OAI221_X1 port map( B1 => n13712, B2 => n16888, C1 => n13424, C2 =>
                           n16885, A => n15594, ZN => n15590);
   U15038 : AOI22_X1 port map( A1 => n16882, A2 => n14923, B1 => n16880, B2 => 
                           n14947, ZN => n15594);
   U15039 : OAI221_X1 port map( B1 => n13711, B2 => n16888, C1 => n13423, C2 =>
                           n16885, A => n15577, ZN => n15573);
   U15040 : AOI22_X1 port map( A1 => n16882, A2 => n14922, B1 => n16880, B2 => 
                           n14946, ZN => n15577);
   U15041 : OAI221_X1 port map( B1 => n13710, B2 => n16888, C1 => n13422, C2 =>
                           n16885, A => n15560, ZN => n15556);
   U15042 : AOI22_X1 port map( A1 => n16882, A2 => n14921, B1 => n16880, B2 => 
                           n14945, ZN => n15560);
   U15043 : OAI221_X1 port map( B1 => n13709, B2 => n16889, C1 => n13421, C2 =>
                           n16886, A => n15543, ZN => n15539);
   U15044 : AOI22_X1 port map( A1 => n16883, A2 => n14920, B1 => n16880, B2 => 
                           n14944, ZN => n15543);
   U15045 : OAI221_X1 port map( B1 => n13708, B2 => n16889, C1 => n13420, C2 =>
                           n16886, A => n15526, ZN => n15522);
   U15046 : AOI22_X1 port map( A1 => n16883, A2 => n14919, B1 => n16880, B2 => 
                           n14943, ZN => n15526);
   U15047 : OAI221_X1 port map( B1 => n13707, B2 => n16889, C1 => n13419, C2 =>
                           n16886, A => n15509, ZN => n15505);
   U15048 : AOI22_X1 port map( A1 => n16883, A2 => n14918, B1 => n16880, B2 => 
                           n14942, ZN => n15509);
   U15049 : OAI221_X1 port map( B1 => n13706, B2 => n16889, C1 => n13418, C2 =>
                           n16886, A => n15492, ZN => n15488);
   U15050 : AOI22_X1 port map( A1 => n16883, A2 => n14917, B1 => n16880, B2 => 
                           n14941, ZN => n15492);
   U15051 : OAI221_X1 port map( B1 => n13705, B2 => n16889, C1 => n13417, C2 =>
                           n16886, A => n15475, ZN => n15471);
   U15052 : AOI22_X1 port map( A1 => n16883, A2 => n14916, B1 => n16880, B2 => 
                           n14940, ZN => n15475);
   U15053 : OAI221_X1 port map( B1 => n13704, B2 => n16889, C1 => n13416, C2 =>
                           n16886, A => n15458, ZN => n15454);
   U15054 : AOI22_X1 port map( A1 => n16883, A2 => n14915, B1 => n16880, B2 => 
                           n14939, ZN => n15458);
   U15055 : OAI221_X1 port map( B1 => n13703, B2 => n16889, C1 => n13415, C2 =>
                           n16886, A => n15441, ZN => n15437);
   U15056 : AOI22_X1 port map( A1 => n16883, A2 => n14914, B1 => n16880, B2 => 
                           n14938, ZN => n15441);
   U15057 : OAI221_X1 port map( B1 => n13702, B2 => n16889, C1 => n13414, C2 =>
                           n16886, A => n15424, ZN => n15420);
   U15058 : AOI22_X1 port map( A1 => n16883, A2 => n14913, B1 => n16880, B2 => 
                           n14937, ZN => n15424);
   U15059 : OAI221_X1 port map( B1 => n13701, B2 => n16889, C1 => n13413, C2 =>
                           n16886, A => n15407, ZN => n15403);
   U15060 : AOI22_X1 port map( A1 => n16883, A2 => n14912, B1 => n16879, B2 => 
                           n14936, ZN => n15407);
   U15061 : OAI221_X1 port map( B1 => n13700, B2 => n16889, C1 => n13412, C2 =>
                           n16886, A => n15390, ZN => n15386);
   U15062 : AOI22_X1 port map( A1 => n16883, A2 => n14911, B1 => n16879, B2 => 
                           n14935, ZN => n15390);
   U15063 : OAI221_X1 port map( B1 => n13699, B2 => n16889, C1 => n13411, C2 =>
                           n16886, A => n15373, ZN => n15369);
   U15064 : AOI22_X1 port map( A1 => n16883, A2 => n14910, B1 => n16879, B2 => 
                           n14934, ZN => n15373);
   U15065 : OAI221_X1 port map( B1 => n13698, B2 => n16889, C1 => n13410, C2 =>
                           n16886, A => n15356, ZN => n15352);
   U15066 : AOI22_X1 port map( A1 => n16883, A2 => n14909, B1 => n16879, B2 => 
                           n14933, ZN => n15356);
   U15067 : OAI221_X1 port map( B1 => n13529, B2 => n16774, C1 => n13593, C2 =>
                           n16771, A => n16336, ZN => n16333);
   U15068 : AOI22_X1 port map( A1 => n16768, A2 => n14980, B1 => n16767, B2 => 
                           n15004, ZN => n16336);
   U15069 : OAI221_X1 port map( B1 => n13520, B2 => n16774, C1 => n13584, C2 =>
                           n16771, A => n16178, ZN => n16176);
   U15070 : AOI22_X1 port map( A1 => n16768, A2 => n14971, B1 => n16766, B2 => 
                           n14995, ZN => n16178);
   U15071 : OAI221_X1 port map( B1 => n13519, B2 => n16774, C1 => n13583, C2 =>
                           n16771, A => n16161, ZN => n16159);
   U15072 : AOI22_X1 port map( A1 => n16768, A2 => n14970, B1 => n16766, B2 => 
                           n14994, ZN => n16161);
   U15073 : OAI221_X1 port map( B1 => n13518, B2 => n16774, C1 => n13582, C2 =>
                           n16771, A => n16144, ZN => n16142);
   U15074 : AOI22_X1 port map( A1 => n16768, A2 => n14969, B1 => n16766, B2 => 
                           n14993, ZN => n16144);
   U15075 : OAI221_X1 port map( B1 => n13517, B2 => n16775, C1 => n13581, C2 =>
                           n16772, A => n16127, ZN => n16125);
   U15076 : AOI22_X1 port map( A1 => n16769, A2 => n14968, B1 => n16766, B2 => 
                           n14992, ZN => n16127);
   U15077 : OAI221_X1 port map( B1 => n13516, B2 => n16775, C1 => n13580, C2 =>
                           n16772, A => n16110, ZN => n16108);
   U15078 : AOI22_X1 port map( A1 => n16769, A2 => n14967, B1 => n16766, B2 => 
                           n14991, ZN => n16110);
   U15079 : OAI221_X1 port map( B1 => n13515, B2 => n16775, C1 => n13579, C2 =>
                           n16772, A => n16093, ZN => n16091);
   U15080 : AOI22_X1 port map( A1 => n16769, A2 => n14966, B1 => n16766, B2 => 
                           n14990, ZN => n16093);
   U15081 : OAI221_X1 port map( B1 => n13514, B2 => n16775, C1 => n13578, C2 =>
                           n16772, A => n16076, ZN => n16074);
   U15082 : AOI22_X1 port map( A1 => n16769, A2 => n14965, B1 => n16766, B2 => 
                           n14989, ZN => n16076);
   U15083 : OAI221_X1 port map( B1 => n13513, B2 => n16775, C1 => n13577, C2 =>
                           n16772, A => n16059, ZN => n16057);
   U15084 : AOI22_X1 port map( A1 => n16769, A2 => n14964, B1 => n16766, B2 => 
                           n14988, ZN => n16059);
   U15085 : OAI221_X1 port map( B1 => n13512, B2 => n16775, C1 => n13576, C2 =>
                           n16772, A => n16042, ZN => n16040);
   U15086 : AOI22_X1 port map( A1 => n16769, A2 => n14963, B1 => n16766, B2 => 
                           n14987, ZN => n16042);
   U15087 : OAI221_X1 port map( B1 => n13511, B2 => n16775, C1 => n13575, C2 =>
                           n16772, A => n16025, ZN => n16023);
   U15088 : AOI22_X1 port map( A1 => n16769, A2 => n14962, B1 => n16766, B2 => 
                           n14986, ZN => n16025);
   U15089 : OAI221_X1 port map( B1 => n13510, B2 => n16775, C1 => n13574, C2 =>
                           n16772, A => n16008, ZN => n16006);
   U15090 : AOI22_X1 port map( A1 => n16769, A2 => n14961, B1 => n16766, B2 => 
                           n14985, ZN => n16008);
   U15091 : OAI221_X1 port map( B1 => n13509, B2 => n16775, C1 => n13573, C2 =>
                           n16772, A => n15991, ZN => n15989);
   U15092 : AOI22_X1 port map( A1 => n16769, A2 => n14960, B1 => n16765, B2 => 
                           n14984, ZN => n15991);
   U15093 : OAI221_X1 port map( B1 => n13508, B2 => n16775, C1 => n13572, C2 =>
                           n16772, A => n15974, ZN => n15972);
   U15094 : AOI22_X1 port map( A1 => n16769, A2 => n14959, B1 => n16765, B2 => 
                           n14983, ZN => n15974);
   U15095 : OAI221_X1 port map( B1 => n13507, B2 => n16775, C1 => n13571, C2 =>
                           n16772, A => n15957, ZN => n15955);
   U15096 : AOI22_X1 port map( A1 => n16769, A2 => n14958, B1 => n16765, B2 => 
                           n14982, ZN => n15957);
   U15097 : OAI221_X1 port map( B1 => n13506, B2 => n16775, C1 => n13570, C2 =>
                           n16772, A => n15940, ZN => n15938);
   U15098 : AOI22_X1 port map( A1 => n16769, A2 => n14957, B1 => n16765, B2 => 
                           n14981, ZN => n15940);
   U15099 : OAI221_X1 port map( B1 => n13529, B2 => n16867, C1 => n13593, C2 =>
                           n16864, A => n15755, ZN => n15752);
   U15100 : AOI22_X1 port map( A1 => n16861, A2 => n14980, B1 => n16860, B2 => 
                           n15004, ZN => n15755);
   U15101 : OAI221_X1 port map( B1 => n13520, B2 => n16867, C1 => n13584, C2 =>
                           n16864, A => n15597, ZN => n15595);
   U15102 : AOI22_X1 port map( A1 => n16861, A2 => n14971, B1 => n16859, B2 => 
                           n14995, ZN => n15597);
   U15103 : OAI221_X1 port map( B1 => n13519, B2 => n16867, C1 => n13583, C2 =>
                           n16864, A => n15580, ZN => n15578);
   U15104 : AOI22_X1 port map( A1 => n16861, A2 => n14970, B1 => n16859, B2 => 
                           n14994, ZN => n15580);
   U15105 : OAI221_X1 port map( B1 => n13518, B2 => n16867, C1 => n13582, C2 =>
                           n16864, A => n15563, ZN => n15561);
   U15106 : AOI22_X1 port map( A1 => n16861, A2 => n14969, B1 => n16859, B2 => 
                           n14993, ZN => n15563);
   U15107 : OAI221_X1 port map( B1 => n13517, B2 => n16868, C1 => n13581, C2 =>
                           n16865, A => n15546, ZN => n15544);
   U15108 : AOI22_X1 port map( A1 => n16862, A2 => n14968, B1 => n16859, B2 => 
                           n14992, ZN => n15546);
   U15109 : OAI221_X1 port map( B1 => n13516, B2 => n16868, C1 => n13580, C2 =>
                           n16865, A => n15529, ZN => n15527);
   U15110 : AOI22_X1 port map( A1 => n16862, A2 => n14967, B1 => n16859, B2 => 
                           n14991, ZN => n15529);
   U15111 : OAI221_X1 port map( B1 => n13515, B2 => n16868, C1 => n13579, C2 =>
                           n16865, A => n15512, ZN => n15510);
   U15112 : AOI22_X1 port map( A1 => n16862, A2 => n14966, B1 => n16859, B2 => 
                           n14990, ZN => n15512);
   U15113 : OAI221_X1 port map( B1 => n13514, B2 => n16868, C1 => n13578, C2 =>
                           n16865, A => n15495, ZN => n15493);
   U15114 : AOI22_X1 port map( A1 => n16862, A2 => n14965, B1 => n16859, B2 => 
                           n14989, ZN => n15495);
   U15115 : OAI221_X1 port map( B1 => n13513, B2 => n16868, C1 => n13577, C2 =>
                           n16865, A => n15478, ZN => n15476);
   U15116 : AOI22_X1 port map( A1 => n16862, A2 => n14964, B1 => n16859, B2 => 
                           n14988, ZN => n15478);
   U15117 : OAI221_X1 port map( B1 => n13512, B2 => n16868, C1 => n13576, C2 =>
                           n16865, A => n15461, ZN => n15459);
   U15118 : AOI22_X1 port map( A1 => n16862, A2 => n14963, B1 => n16859, B2 => 
                           n14987, ZN => n15461);
   U15119 : OAI221_X1 port map( B1 => n13511, B2 => n16868, C1 => n13575, C2 =>
                           n16865, A => n15444, ZN => n15442);
   U15120 : AOI22_X1 port map( A1 => n16862, A2 => n14962, B1 => n16859, B2 => 
                           n14986, ZN => n15444);
   U15121 : OAI221_X1 port map( B1 => n13510, B2 => n16868, C1 => n13574, C2 =>
                           n16865, A => n15427, ZN => n15425);
   U15122 : AOI22_X1 port map( A1 => n16862, A2 => n14961, B1 => n16859, B2 => 
                           n14985, ZN => n15427);
   U15123 : OAI221_X1 port map( B1 => n13509, B2 => n16868, C1 => n13573, C2 =>
                           n16865, A => n15410, ZN => n15408);
   U15124 : AOI22_X1 port map( A1 => n16862, A2 => n14960, B1 => n16858, B2 => 
                           n14984, ZN => n15410);
   U15125 : OAI221_X1 port map( B1 => n13508, B2 => n16868, C1 => n13572, C2 =>
                           n16865, A => n15393, ZN => n15391);
   U15126 : AOI22_X1 port map( A1 => n16862, A2 => n14959, B1 => n16858, B2 => 
                           n14983, ZN => n15393);
   U15127 : OAI221_X1 port map( B1 => n13507, B2 => n16868, C1 => n13571, C2 =>
                           n16865, A => n15376, ZN => n15374);
   U15128 : AOI22_X1 port map( A1 => n16862, A2 => n14958, B1 => n16858, B2 => 
                           n14982, ZN => n15376);
   U15129 : OAI221_X1 port map( B1 => n13506, B2 => n16868, C1 => n13570, C2 =>
                           n16865, A => n15359, ZN => n15357);
   U15130 : AOI22_X1 port map( A1 => n16862, A2 => n14957, B1 => n16858, B2 => 
                           n14981, ZN => n15359);
   U15131 : OAI22_X1 port map( A1 => n13473, A2 => n16740, B1 => n13729, B2 => 
                           n16739, ZN => n15927);
   U15132 : OAI22_X1 port map( A1 => n13472, A2 => n16741, B1 => n13728, B2 => 
                           n16739, ZN => n15910);
   U15133 : OAI22_X1 port map( A1 => n13471, A2 => n16740, B1 => n13727, B2 => 
                           n16739, ZN => n15893);
   U15134 : OAI22_X1 port map( A1 => n13470, A2 => n16741, B1 => n13726, B2 => 
                           n16739, ZN => n15876);
   U15135 : OAI22_X1 port map( A1 => n13469, A2 => n16740, B1 => n13725, B2 => 
                           n16739, ZN => n15859);
   U15136 : OAI22_X1 port map( A1 => n13468, A2 => n16741, B1 => n13724, B2 => 
                           n16739, ZN => n15842);
   U15137 : OAI22_X1 port map( A1 => n13467, A2 => n16740, B1 => n13723, B2 => 
                           n16739, ZN => n15825);
   U15138 : OAI22_X1 port map( A1 => n13466, A2 => n16741, B1 => n13722, B2 => 
                           n16739, ZN => n15804);
   U15139 : OAI22_X1 port map( A1 => n13473, A2 => n16833, B1 => n13729, B2 => 
                           n16832, ZN => n15346);
   U15140 : OAI22_X1 port map( A1 => n13472, A2 => n16834, B1 => n13728, B2 => 
                           n16832, ZN => n15329);
   U15141 : OAI22_X1 port map( A1 => n13471, A2 => n16833, B1 => n13727, B2 => 
                           n16832, ZN => n15312);
   U15142 : OAI22_X1 port map( A1 => n13470, A2 => n16834, B1 => n13726, B2 => 
                           n16832, ZN => n15295);
   U15143 : OAI22_X1 port map( A1 => n13469, A2 => n16833, B1 => n13725, B2 => 
                           n16832, ZN => n15278);
   U15144 : OAI22_X1 port map( A1 => n13468, A2 => n16834, B1 => n13724, B2 => 
                           n16832, ZN => n15261);
   U15145 : OAI22_X1 port map( A1 => n13467, A2 => n16833, B1 => n13723, B2 => 
                           n16832, ZN => n15244);
   U15146 : OAI22_X1 port map( A1 => n13466, A2 => n16834, B1 => n13722, B2 => 
                           n16832, ZN => n15223);
   U15147 : OAI22_X1 port map( A1 => n13345, A2 => n17308, B1 => n13601, B2 => 
                           n17305, ZN => n15928);
   U15148 : OAI22_X1 port map( A1 => n13344, A2 => n17308, B1 => n13600, B2 => 
                           n17305, ZN => n15911);
   U15149 : OAI22_X1 port map( A1 => n13343, A2 => n17308, B1 => n13599, B2 => 
                           n17305, ZN => n15894);
   U15150 : OAI22_X1 port map( A1 => n13342, A2 => n17308, B1 => n13598, B2 => 
                           n17305, ZN => n15877);
   U15151 : OAI22_X1 port map( A1 => n13341, A2 => n17308, B1 => n13597, B2 => 
                           n17305, ZN => n15860);
   U15152 : OAI22_X1 port map( A1 => n13340, A2 => n17308, B1 => n13596, B2 => 
                           n17305, ZN => n15843);
   U15153 : OAI22_X1 port map( A1 => n13339, A2 => n17308, B1 => n13595, B2 => 
                           n17305, ZN => n15826);
   U15154 : OAI22_X1 port map( A1 => n13338, A2 => n17308, B1 => n13594, B2 => 
                           n17305, ZN => n15809);
   U15155 : OAI22_X1 port map( A1 => n13345, A2 => n17314, B1 => n13601, B2 => 
                           n17311, ZN => n15347);
   U15156 : OAI22_X1 port map( A1 => n13344, A2 => n17314, B1 => n13600, B2 => 
                           n17311, ZN => n15330);
   U15157 : OAI22_X1 port map( A1 => n13343, A2 => n17314, B1 => n13599, B2 => 
                           n17311, ZN => n15313);
   U15158 : OAI22_X1 port map( A1 => n13342, A2 => n17314, B1 => n13598, B2 => 
                           n17311, ZN => n15296);
   U15159 : OAI22_X1 port map( A1 => n13341, A2 => n17314, B1 => n13597, B2 => 
                           n17311, ZN => n15279);
   U15160 : OAI22_X1 port map( A1 => n13340, A2 => n17314, B1 => n13596, B2 => 
                           n17311, ZN => n15262);
   U15161 : OAI22_X1 port map( A1 => n13339, A2 => n17314, B1 => n13595, B2 => 
                           n17311, ZN => n15245);
   U15162 : OAI22_X1 port map( A1 => n13338, A2 => n17314, B1 => n13594, B2 => 
                           n17311, ZN => n15228);
   U15163 : OAI22_X1 port map( A1 => n13497, A2 => n16740, B1 => n13753, B2 => 
                           n16738, ZN => n16340);
   U15164 : OAI22_X1 port map( A1 => n13496, A2 => n16740, B1 => n13752, B2 => 
                           n16738, ZN => n16318);
   U15165 : OAI22_X1 port map( A1 => n13495, A2 => n16740, B1 => n13751, B2 => 
                           n16738, ZN => n16301);
   U15166 : OAI22_X1 port map( A1 => n13494, A2 => n16740, B1 => n13750, B2 => 
                           n16738, ZN => n16284);
   U15167 : OAI22_X1 port map( A1 => n13493, A2 => n16740, B1 => n13749, B2 => 
                           n16738, ZN => n16267);
   U15168 : OAI22_X1 port map( A1 => n13492, A2 => n16740, B1 => n13748, B2 => 
                           n16738, ZN => n16250);
   U15169 : OAI22_X1 port map( A1 => n13491, A2 => n16740, B1 => n13747, B2 => 
                           n16738, ZN => n16233);
   U15170 : OAI22_X1 port map( A1 => n13490, A2 => n16740, B1 => n13746, B2 => 
                           n16738, ZN => n16216);
   U15171 : OAI22_X1 port map( A1 => n13489, A2 => n16740, B1 => n13745, B2 => 
                           n16738, ZN => n16199);
   U15172 : OAI22_X1 port map( A1 => n13488, A2 => n16740, B1 => n13744, B2 => 
                           n16738, ZN => n16182);
   U15173 : OAI22_X1 port map( A1 => n13487, A2 => n16740, B1 => n13743, B2 => 
                           n16738, ZN => n16165);
   U15174 : OAI22_X1 port map( A1 => n13486, A2 => n16740, B1 => n13742, B2 => 
                           n16738, ZN => n16148);
   U15175 : OAI22_X1 port map( A1 => n13485, A2 => n16741, B1 => n13741, B2 => 
                           n16739, ZN => n16131);
   U15176 : OAI22_X1 port map( A1 => n13484, A2 => n16741, B1 => n13740, B2 => 
                           n16739, ZN => n16114);
   U15177 : OAI22_X1 port map( A1 => n13483, A2 => n16741, B1 => n13739, B2 => 
                           n16739, ZN => n16097);
   U15178 : OAI22_X1 port map( A1 => n13482, A2 => n16741, B1 => n13738, B2 => 
                           n16739, ZN => n16080);
   U15179 : OAI22_X1 port map( A1 => n13481, A2 => n16741, B1 => n13737, B2 => 
                           n16738, ZN => n16063);
   U15180 : OAI22_X1 port map( A1 => n13480, A2 => n16741, B1 => n13736, B2 => 
                           n16739, ZN => n16046);
   U15181 : OAI22_X1 port map( A1 => n13479, A2 => n16741, B1 => n13735, B2 => 
                           n16738, ZN => n16029);
   U15182 : OAI22_X1 port map( A1 => n13478, A2 => n16741, B1 => n13734, B2 => 
                           n16739, ZN => n16012);
   U15183 : OAI22_X1 port map( A1 => n13477, A2 => n16741, B1 => n13733, B2 => 
                           n16738, ZN => n15995);
   U15184 : OAI22_X1 port map( A1 => n13476, A2 => n16741, B1 => n13732, B2 => 
                           n16739, ZN => n15978);
   U15185 : OAI22_X1 port map( A1 => n13475, A2 => n16741, B1 => n13731, B2 => 
                           n16738, ZN => n15961);
   U15186 : OAI22_X1 port map( A1 => n13474, A2 => n16741, B1 => n13730, B2 => 
                           n16739, ZN => n15944);
   U15187 : OAI22_X1 port map( A1 => n13497, A2 => n16833, B1 => n13753, B2 => 
                           n16831, ZN => n15759);
   U15188 : OAI22_X1 port map( A1 => n13496, A2 => n16833, B1 => n13752, B2 => 
                           n16831, ZN => n15737);
   U15189 : OAI22_X1 port map( A1 => n13495, A2 => n16833, B1 => n13751, B2 => 
                           n16831, ZN => n15720);
   U15190 : OAI22_X1 port map( A1 => n13494, A2 => n16833, B1 => n13750, B2 => 
                           n16831, ZN => n15703);
   U15191 : OAI22_X1 port map( A1 => n13493, A2 => n16833, B1 => n13749, B2 => 
                           n16831, ZN => n15686);
   U15192 : OAI22_X1 port map( A1 => n13492, A2 => n16833, B1 => n13748, B2 => 
                           n16831, ZN => n15669);
   U15193 : OAI22_X1 port map( A1 => n13491, A2 => n16833, B1 => n13747, B2 => 
                           n16831, ZN => n15652);
   U15194 : OAI22_X1 port map( A1 => n13490, A2 => n16833, B1 => n13746, B2 => 
                           n16831, ZN => n15635);
   U15195 : OAI22_X1 port map( A1 => n13489, A2 => n16833, B1 => n13745, B2 => 
                           n16831, ZN => n15618);
   U15196 : OAI22_X1 port map( A1 => n13488, A2 => n16833, B1 => n13744, B2 => 
                           n16831, ZN => n15601);
   U15197 : OAI22_X1 port map( A1 => n13487, A2 => n16833, B1 => n13743, B2 => 
                           n16831, ZN => n15584);
   U15198 : OAI22_X1 port map( A1 => n13486, A2 => n16833, B1 => n13742, B2 => 
                           n16831, ZN => n15567);
   U15199 : OAI22_X1 port map( A1 => n13485, A2 => n16834, B1 => n13741, B2 => 
                           n16832, ZN => n15550);
   U15200 : OAI22_X1 port map( A1 => n13484, A2 => n16834, B1 => n13740, B2 => 
                           n16832, ZN => n15533);
   U15201 : OAI22_X1 port map( A1 => n13483, A2 => n16834, B1 => n13739, B2 => 
                           n16832, ZN => n15516);
   U15202 : OAI22_X1 port map( A1 => n13482, A2 => n16834, B1 => n13738, B2 => 
                           n16832, ZN => n15499);
   U15203 : OAI22_X1 port map( A1 => n13481, A2 => n16834, B1 => n13737, B2 => 
                           n16831, ZN => n15482);
   U15204 : OAI22_X1 port map( A1 => n13480, A2 => n16834, B1 => n13736, B2 => 
                           n16832, ZN => n15465);
   U15205 : OAI22_X1 port map( A1 => n13479, A2 => n16834, B1 => n13735, B2 => 
                           n16831, ZN => n15448);
   U15206 : OAI22_X1 port map( A1 => n13478, A2 => n16834, B1 => n13734, B2 => 
                           n16832, ZN => n15431);
   U15207 : OAI22_X1 port map( A1 => n13477, A2 => n16834, B1 => n13733, B2 => 
                           n16831, ZN => n15414);
   U15208 : OAI22_X1 port map( A1 => n13476, A2 => n16834, B1 => n13732, B2 => 
                           n16832, ZN => n15397);
   U15209 : OAI22_X1 port map( A1 => n13475, A2 => n16834, B1 => n13731, B2 => 
                           n16831, ZN => n15380);
   U15210 : OAI22_X1 port map( A1 => n13474, A2 => n16834, B1 => n13730, B2 => 
                           n16832, ZN => n15363);
   U15211 : OAI22_X1 port map( A1 => n13369, A2 => n17306, B1 => n13625, B2 => 
                           n17303, ZN => n16341);
   U15212 : OAI22_X1 port map( A1 => n13368, A2 => n17306, B1 => n13624, B2 => 
                           n17303, ZN => n16319);
   U15213 : OAI22_X1 port map( A1 => n13367, A2 => n17306, B1 => n13623, B2 => 
                           n17303, ZN => n16302);
   U15214 : OAI22_X1 port map( A1 => n13366, A2 => n17306, B1 => n13622, B2 => 
                           n17303, ZN => n16285);
   U15215 : OAI22_X1 port map( A1 => n13365, A2 => n17306, B1 => n13621, B2 => 
                           n17303, ZN => n16268);
   U15216 : OAI22_X1 port map( A1 => n13364, A2 => n17306, B1 => n13620, B2 => 
                           n17303, ZN => n16251);
   U15217 : OAI22_X1 port map( A1 => n13363, A2 => n17306, B1 => n13619, B2 => 
                           n17303, ZN => n16234);
   U15218 : OAI22_X1 port map( A1 => n13362, A2 => n17306, B1 => n13618, B2 => 
                           n17303, ZN => n16217);
   U15219 : OAI22_X1 port map( A1 => n13361, A2 => n17306, B1 => n13617, B2 => 
                           n17303, ZN => n16200);
   U15220 : OAI22_X1 port map( A1 => n13360, A2 => n17306, B1 => n13616, B2 => 
                           n17303, ZN => n16183);
   U15221 : OAI22_X1 port map( A1 => n13359, A2 => n17306, B1 => n13615, B2 => 
                           n17303, ZN => n16166);
   U15222 : OAI22_X1 port map( A1 => n13358, A2 => n17306, B1 => n13614, B2 => 
                           n17303, ZN => n16149);
   U15223 : OAI22_X1 port map( A1 => n13357, A2 => n17307, B1 => n13613, B2 => 
                           n17304, ZN => n16132);
   U15224 : OAI22_X1 port map( A1 => n13356, A2 => n17307, B1 => n13612, B2 => 
                           n17304, ZN => n16115);
   U15225 : OAI22_X1 port map( A1 => n13355, A2 => n17307, B1 => n13611, B2 => 
                           n17304, ZN => n16098);
   U15226 : OAI22_X1 port map( A1 => n13354, A2 => n17307, B1 => n13610, B2 => 
                           n17304, ZN => n16081);
   U15227 : OAI22_X1 port map( A1 => n13353, A2 => n17307, B1 => n13609, B2 => 
                           n17304, ZN => n16064);
   U15228 : OAI22_X1 port map( A1 => n13352, A2 => n17307, B1 => n13608, B2 => 
                           n17304, ZN => n16047);
   U15229 : OAI22_X1 port map( A1 => n13351, A2 => n17307, B1 => n13607, B2 => 
                           n17304, ZN => n16030);
   U15230 : OAI22_X1 port map( A1 => n13350, A2 => n17307, B1 => n13606, B2 => 
                           n17304, ZN => n16013);
   U15231 : OAI22_X1 port map( A1 => n13349, A2 => n17307, B1 => n13605, B2 => 
                           n17304, ZN => n15996);
   U15232 : OAI22_X1 port map( A1 => n13348, A2 => n17307, B1 => n13604, B2 => 
                           n17304, ZN => n15979);
   U15233 : OAI22_X1 port map( A1 => n13347, A2 => n17307, B1 => n13603, B2 => 
                           n17304, ZN => n15962);
   U15234 : OAI22_X1 port map( A1 => n13346, A2 => n17307, B1 => n13602, B2 => 
                           n17304, ZN => n15945);
   U15235 : OAI22_X1 port map( A1 => n13369, A2 => n17312, B1 => n13625, B2 => 
                           n17309, ZN => n15760);
   U15236 : OAI22_X1 port map( A1 => n13368, A2 => n17312, B1 => n13624, B2 => 
                           n17309, ZN => n15738);
   U15237 : OAI22_X1 port map( A1 => n13367, A2 => n17312, B1 => n13623, B2 => 
                           n17309, ZN => n15721);
   U15238 : OAI22_X1 port map( A1 => n13366, A2 => n17312, B1 => n13622, B2 => 
                           n17309, ZN => n15704);
   U15239 : OAI22_X1 port map( A1 => n13365, A2 => n17312, B1 => n13621, B2 => 
                           n17309, ZN => n15687);
   U15240 : OAI22_X1 port map( A1 => n13364, A2 => n17312, B1 => n13620, B2 => 
                           n17309, ZN => n15670);
   U15241 : OAI22_X1 port map( A1 => n13363, A2 => n17312, B1 => n13619, B2 => 
                           n17309, ZN => n15653);
   U15242 : OAI22_X1 port map( A1 => n13362, A2 => n17312, B1 => n13618, B2 => 
                           n17309, ZN => n15636);
   U15243 : OAI22_X1 port map( A1 => n13361, A2 => n17312, B1 => n13617, B2 => 
                           n17309, ZN => n15619);
   U15244 : OAI22_X1 port map( A1 => n13360, A2 => n17312, B1 => n13616, B2 => 
                           n17309, ZN => n15602);
   U15245 : OAI22_X1 port map( A1 => n13359, A2 => n17312, B1 => n13615, B2 => 
                           n17309, ZN => n15585);
   U15246 : OAI22_X1 port map( A1 => n13358, A2 => n17312, B1 => n13614, B2 => 
                           n17309, ZN => n15568);
   U15247 : OAI22_X1 port map( A1 => n13357, A2 => n17313, B1 => n13613, B2 => 
                           n17310, ZN => n15551);
   U15248 : OAI22_X1 port map( A1 => n13356, A2 => n17313, B1 => n13612, B2 => 
                           n17310, ZN => n15534);
   U15249 : OAI22_X1 port map( A1 => n13355, A2 => n17313, B1 => n13611, B2 => 
                           n17310, ZN => n15517);
   U15250 : OAI22_X1 port map( A1 => n13354, A2 => n17313, B1 => n13610, B2 => 
                           n17310, ZN => n15500);
   U15251 : OAI22_X1 port map( A1 => n13353, A2 => n17313, B1 => n13609, B2 => 
                           n17310, ZN => n15483);
   U15252 : OAI22_X1 port map( A1 => n13352, A2 => n17313, B1 => n13608, B2 => 
                           n17310, ZN => n15466);
   U15253 : OAI22_X1 port map( A1 => n13351, A2 => n17313, B1 => n13607, B2 => 
                           n17310, ZN => n15449);
   U15254 : OAI22_X1 port map( A1 => n13350, A2 => n17313, B1 => n13606, B2 => 
                           n17310, ZN => n15432);
   U15255 : OAI22_X1 port map( A1 => n13349, A2 => n17313, B1 => n13605, B2 => 
                           n17310, ZN => n15415);
   U15256 : OAI22_X1 port map( A1 => n13348, A2 => n17313, B1 => n13604, B2 => 
                           n17310, ZN => n15398);
   U15257 : OAI22_X1 port map( A1 => n13347, A2 => n17313, B1 => n13603, B2 => 
                           n17310, ZN => n15381);
   U15258 : OAI22_X1 port map( A1 => n13346, A2 => n17313, B1 => n13602, B2 => 
                           n17310, ZN => n15364);
   U15259 : OAI22_X1 port map( A1 => n14693, A2 => n16782, B1 => n13313, B2 => 
                           n16779, ZN => n15922);
   U15260 : OAI22_X1 port map( A1 => n14692, A2 => n16782, B1 => n13312, B2 => 
                           n16779, ZN => n15905);
   U15261 : OAI22_X1 port map( A1 => n14691, A2 => n16782, B1 => n13311, B2 => 
                           n16779, ZN => n15888);
   U15262 : OAI22_X1 port map( A1 => n14690, A2 => n16782, B1 => n13310, B2 => 
                           n16779, ZN => n15871);
   U15263 : OAI22_X1 port map( A1 => n14689, A2 => n16782, B1 => n13309, B2 => 
                           n16779, ZN => n15854);
   U15264 : OAI22_X1 port map( A1 => n14688, A2 => n16782, B1 => n13308, B2 => 
                           n16779, ZN => n15837);
   U15265 : OAI22_X1 port map( A1 => n14687, A2 => n16782, B1 => n13307, B2 => 
                           n16779, ZN => n15820);
   U15266 : OAI22_X1 port map( A1 => n14686, A2 => n16782, B1 => n13306, B2 => 
                           n16779, ZN => n15785);
   U15267 : OAI22_X1 port map( A1 => n14693, A2 => n16875, B1 => n13313, B2 => 
                           n16872, ZN => n15341);
   U15268 : OAI22_X1 port map( A1 => n14692, A2 => n16875, B1 => n13312, B2 => 
                           n16872, ZN => n15324);
   U15269 : OAI22_X1 port map( A1 => n14691, A2 => n16875, B1 => n13311, B2 => 
                           n16872, ZN => n15307);
   U15270 : OAI22_X1 port map( A1 => n14690, A2 => n16875, B1 => n13310, B2 => 
                           n16872, ZN => n15290);
   U15271 : OAI22_X1 port map( A1 => n14689, A2 => n16875, B1 => n13309, B2 => 
                           n16872, ZN => n15273);
   U15272 : OAI22_X1 port map( A1 => n14688, A2 => n16875, B1 => n13308, B2 => 
                           n16872, ZN => n15256);
   U15273 : OAI22_X1 port map( A1 => n14687, A2 => n16875, B1 => n13307, B2 => 
                           n16872, ZN => n15239);
   U15274 : OAI22_X1 port map( A1 => n14686, A2 => n16875, B1 => n13306, B2 => 
                           n16872, ZN => n15204);
   U15275 : OAI22_X1 port map( A1 => n14717, A2 => n16780, B1 => n13337, B2 => 
                           n16777, ZN => n16334);
   U15276 : OAI22_X1 port map( A1 => n14716, A2 => n16780, B1 => n13336, B2 => 
                           n16777, ZN => n16313);
   U15277 : OAI22_X1 port map( A1 => n14715, A2 => n16780, B1 => n13335, B2 => 
                           n16777, ZN => n16296);
   U15278 : OAI22_X1 port map( A1 => n14714, A2 => n16780, B1 => n13334, B2 => 
                           n16777, ZN => n16279);
   U15279 : OAI22_X1 port map( A1 => n14713, A2 => n16780, B1 => n13333, B2 => 
                           n16777, ZN => n16262);
   U15280 : OAI22_X1 port map( A1 => n14712, A2 => n16780, B1 => n13332, B2 => 
                           n16777, ZN => n16245);
   U15281 : OAI22_X1 port map( A1 => n14711, A2 => n16780, B1 => n13331, B2 => 
                           n16777, ZN => n16228);
   U15282 : OAI22_X1 port map( A1 => n14710, A2 => n16780, B1 => n13330, B2 => 
                           n16777, ZN => n16211);
   U15283 : OAI22_X1 port map( A1 => n14709, A2 => n16780, B1 => n13329, B2 => 
                           n16777, ZN => n16194);
   U15284 : OAI22_X1 port map( A1 => n14708, A2 => n16780, B1 => n13328, B2 => 
                           n16777, ZN => n16177);
   U15285 : OAI22_X1 port map( A1 => n14707, A2 => n16780, B1 => n13327, B2 => 
                           n16777, ZN => n16160);
   U15286 : OAI22_X1 port map( A1 => n14706, A2 => n16780, B1 => n13326, B2 => 
                           n16777, ZN => n16143);
   U15287 : OAI22_X1 port map( A1 => n14705, A2 => n16781, B1 => n13325, B2 => 
                           n16778, ZN => n16126);
   U15288 : OAI22_X1 port map( A1 => n14704, A2 => n16781, B1 => n13324, B2 => 
                           n16778, ZN => n16109);
   U15289 : OAI22_X1 port map( A1 => n14703, A2 => n16781, B1 => n13323, B2 => 
                           n16778, ZN => n16092);
   U15290 : OAI22_X1 port map( A1 => n14702, A2 => n16781, B1 => n13322, B2 => 
                           n16778, ZN => n16075);
   U15291 : OAI22_X1 port map( A1 => n14701, A2 => n16781, B1 => n13321, B2 => 
                           n16778, ZN => n16058);
   U15292 : OAI22_X1 port map( A1 => n14700, A2 => n16781, B1 => n13320, B2 => 
                           n16778, ZN => n16041);
   U15293 : OAI22_X1 port map( A1 => n14699, A2 => n16781, B1 => n13319, B2 => 
                           n16778, ZN => n16024);
   U15294 : OAI22_X1 port map( A1 => n14698, A2 => n16781, B1 => n13318, B2 => 
                           n16778, ZN => n16007);
   U15295 : OAI22_X1 port map( A1 => n14697, A2 => n16781, B1 => n13317, B2 => 
                           n16778, ZN => n15990);
   U15296 : OAI22_X1 port map( A1 => n14696, A2 => n16781, B1 => n13316, B2 => 
                           n16778, ZN => n15973);
   U15297 : OAI22_X1 port map( A1 => n14695, A2 => n16781, B1 => n13315, B2 => 
                           n16778, ZN => n15956);
   U15298 : OAI22_X1 port map( A1 => n14694, A2 => n16781, B1 => n13314, B2 => 
                           n16778, ZN => n15939);
   U15299 : OAI22_X1 port map( A1 => n14717, A2 => n16873, B1 => n13337, B2 => 
                           n16870, ZN => n15753);
   U15300 : OAI22_X1 port map( A1 => n14716, A2 => n16873, B1 => n13336, B2 => 
                           n16870, ZN => n15732);
   U15301 : OAI22_X1 port map( A1 => n14715, A2 => n16873, B1 => n13335, B2 => 
                           n16870, ZN => n15715);
   U15302 : OAI22_X1 port map( A1 => n14714, A2 => n16873, B1 => n13334, B2 => 
                           n16870, ZN => n15698);
   U15303 : OAI22_X1 port map( A1 => n14713, A2 => n16873, B1 => n13333, B2 => 
                           n16870, ZN => n15681);
   U15304 : OAI22_X1 port map( A1 => n14712, A2 => n16873, B1 => n13332, B2 => 
                           n16870, ZN => n15664);
   U15305 : OAI22_X1 port map( A1 => n14711, A2 => n16873, B1 => n13331, B2 => 
                           n16870, ZN => n15647);
   U15306 : OAI22_X1 port map( A1 => n14710, A2 => n16873, B1 => n13330, B2 => 
                           n16870, ZN => n15630);
   U15307 : OAI22_X1 port map( A1 => n14709, A2 => n16873, B1 => n13329, B2 => 
                           n16870, ZN => n15613);
   U15308 : OAI22_X1 port map( A1 => n14708, A2 => n16873, B1 => n13328, B2 => 
                           n16870, ZN => n15596);
   U15309 : OAI22_X1 port map( A1 => n14707, A2 => n16873, B1 => n13327, B2 => 
                           n16870, ZN => n15579);
   U15310 : OAI22_X1 port map( A1 => n14706, A2 => n16873, B1 => n13326, B2 => 
                           n16870, ZN => n15562);
   U15311 : OAI22_X1 port map( A1 => n14705, A2 => n16874, B1 => n13325, B2 => 
                           n16871, ZN => n15545);
   U15312 : OAI22_X1 port map( A1 => n14704, A2 => n16874, B1 => n13324, B2 => 
                           n16871, ZN => n15528);
   U15313 : OAI22_X1 port map( A1 => n14703, A2 => n16874, B1 => n13323, B2 => 
                           n16871, ZN => n15511);
   U15314 : OAI22_X1 port map( A1 => n14702, A2 => n16874, B1 => n13322, B2 => 
                           n16871, ZN => n15494);
   U15315 : OAI22_X1 port map( A1 => n14701, A2 => n16874, B1 => n13321, B2 => 
                           n16871, ZN => n15477);
   U15316 : OAI22_X1 port map( A1 => n14700, A2 => n16874, B1 => n13320, B2 => 
                           n16871, ZN => n15460);
   U15317 : OAI22_X1 port map( A1 => n14699, A2 => n16874, B1 => n13319, B2 => 
                           n16871, ZN => n15443);
   U15318 : OAI22_X1 port map( A1 => n14698, A2 => n16874, B1 => n13318, B2 => 
                           n16871, ZN => n15426);
   U15319 : OAI22_X1 port map( A1 => n14697, A2 => n16874, B1 => n13317, B2 => 
                           n16871, ZN => n15409);
   U15320 : OAI22_X1 port map( A1 => n14696, A2 => n16874, B1 => n13316, B2 => 
                           n16871, ZN => n15392);
   U15321 : OAI22_X1 port map( A1 => n14695, A2 => n16874, B1 => n13315, B2 => 
                           n16871, ZN => n15375);
   U15322 : OAI22_X1 port map( A1 => n14694, A2 => n16874, B1 => n13314, B2 => 
                           n16871, ZN => n15358);
   U15323 : OAI22_X1 port map( A1 => n17113, A2 => n17270, B1 => n15152, B2 => 
                           n14725, ZN => n2036);
   U15324 : OAI22_X1 port map( A1 => n17114, A2 => n17273, B1 => n15152, B2 => 
                           n14724, ZN => n2037);
   U15325 : OAI22_X1 port map( A1 => n17114, A2 => n17276, B1 => n15152, B2 => 
                           n14723, ZN => n2038);
   U15326 : OAI22_X1 port map( A1 => n17114, A2 => n17279, B1 => n15152, B2 => 
                           n14722, ZN => n2039);
   U15327 : OAI22_X1 port map( A1 => n17114, A2 => n17282, B1 => n15152, B2 => 
                           n14721, ZN => n2040);
   U15328 : OAI22_X1 port map( A1 => n17114, A2 => n17285, B1 => n15152, B2 => 
                           n14720, ZN => n2041);
   U15329 : OAI22_X1 port map( A1 => n17115, A2 => n17288, B1 => n15152, B2 => 
                           n14719, ZN => n2042);
   U15330 : OAI22_X1 port map( A1 => n17115, A2 => n17300, B1 => n15152, B2 => 
                           n14718, ZN => n2043);
   U15331 : OAI22_X1 port map( A1 => n17131, A2 => n17270, B1 => n15149, B2 => 
                           n14661, ZN => n2100);
   U15332 : OAI22_X1 port map( A1 => n17132, A2 => n17273, B1 => n15149, B2 => 
                           n14660, ZN => n2101);
   U15333 : OAI22_X1 port map( A1 => n17132, A2 => n17276, B1 => n15149, B2 => 
                           n14659, ZN => n2102);
   U15334 : OAI22_X1 port map( A1 => n17132, A2 => n17279, B1 => n15149, B2 => 
                           n14658, ZN => n2103);
   U15335 : OAI22_X1 port map( A1 => n17132, A2 => n17282, B1 => n15149, B2 => 
                           n14657, ZN => n2104);
   U15336 : OAI22_X1 port map( A1 => n17132, A2 => n17285, B1 => n15149, B2 => 
                           n14656, ZN => n2105);
   U15337 : OAI22_X1 port map( A1 => n17133, A2 => n17288, B1 => n15149, B2 => 
                           n14655, ZN => n2106);
   U15338 : OAI22_X1 port map( A1 => n17133, A2 => n17300, B1 => n15149, B2 => 
                           n14654, ZN => n2107);
   U15339 : OAI22_X1 port map( A1 => n17185, A2 => n17270, B1 => n15139, B2 => 
                           n14533, ZN => n2292);
   U15340 : OAI22_X1 port map( A1 => n17186, A2 => n17273, B1 => n15139, B2 => 
                           n14532, ZN => n2293);
   U15341 : OAI22_X1 port map( A1 => n17186, A2 => n17276, B1 => n15139, B2 => 
                           n14531, ZN => n2294);
   U15342 : OAI22_X1 port map( A1 => n17186, A2 => n17279, B1 => n15139, B2 => 
                           n14530, ZN => n2295);
   U15343 : OAI22_X1 port map( A1 => n17186, A2 => n17282, B1 => n15139, B2 => 
                           n14529, ZN => n2296);
   U15344 : OAI22_X1 port map( A1 => n17186, A2 => n17285, B1 => n15139, B2 => 
                           n14528, ZN => n2297);
   U15345 : OAI22_X1 port map( A1 => n17187, A2 => n17288, B1 => n15139, B2 => 
                           n14527, ZN => n2298);
   U15346 : OAI22_X1 port map( A1 => n17187, A2 => n17300, B1 => n15139, B2 => 
                           n14526, ZN => n2299);
   U15347 : OAI22_X1 port map( A1 => n17194, A2 => n17270, B1 => n15137, B2 => 
                           n14501, ZN => n2324);
   U15348 : OAI22_X1 port map( A1 => n17195, A2 => n17273, B1 => n15137, B2 => 
                           n14500, ZN => n2325);
   U15349 : OAI22_X1 port map( A1 => n17195, A2 => n17276, B1 => n15137, B2 => 
                           n14499, ZN => n2326);
   U15350 : OAI22_X1 port map( A1 => n17195, A2 => n17279, B1 => n15137, B2 => 
                           n14498, ZN => n2327);
   U15351 : OAI22_X1 port map( A1 => n17195, A2 => n17282, B1 => n15137, B2 => 
                           n14497, ZN => n2328);
   U15352 : OAI22_X1 port map( A1 => n17195, A2 => n17285, B1 => n15137, B2 => 
                           n14496, ZN => n2329);
   U15353 : OAI22_X1 port map( A1 => n17196, A2 => n17288, B1 => n15137, B2 => 
                           n14495, ZN => n2330);
   U15354 : OAI22_X1 port map( A1 => n17196, A2 => n17300, B1 => n15137, B2 => 
                           n14494, ZN => n2331);
   U15355 : OAI22_X1 port map( A1 => n17296, A2 => n17270, B1 => n15103, B2 => 
                           n14469, ZN => n2356);
   U15356 : OAI22_X1 port map( A1 => n17297, A2 => n17273, B1 => n15103, B2 => 
                           n14468, ZN => n2357);
   U15357 : OAI22_X1 port map( A1 => n17297, A2 => n17276, B1 => n15103, B2 => 
                           n14467, ZN => n2358);
   U15358 : OAI22_X1 port map( A1 => n17297, A2 => n17279, B1 => n15103, B2 => 
                           n14466, ZN => n2359);
   U15359 : OAI22_X1 port map( A1 => n17297, A2 => n17282, B1 => n15103, B2 => 
                           n14465, ZN => n2360);
   U15360 : OAI22_X1 port map( A1 => n17297, A2 => n17285, B1 => n15103, B2 => 
                           n14464, ZN => n2361);
   U15361 : OAI22_X1 port map( A1 => n17298, A2 => n17288, B1 => n15103, B2 => 
                           n14463, ZN => n2362);
   U15362 : OAI22_X1 port map( A1 => n17298, A2 => n17300, B1 => n15103, B2 => 
                           n14462, ZN => n2363);
   U15363 : OAI22_X1 port map( A1 => n17176, A2 => n17270, B1 => n12833, B2 => 
                           n15141, ZN => n2260);
   U15364 : OAI22_X1 port map( A1 => n17177, A2 => n17273, B1 => n12832, B2 => 
                           n15141, ZN => n2261);
   U15365 : OAI22_X1 port map( A1 => n17177, A2 => n17276, B1 => n12831, B2 => 
                           n15141, ZN => n2262);
   U15366 : OAI22_X1 port map( A1 => n17177, A2 => n17279, B1 => n12830, B2 => 
                           n15141, ZN => n2263);
   U15367 : OAI22_X1 port map( A1 => n17177, A2 => n17282, B1 => n12829, B2 => 
                           n15141, ZN => n2264);
   U15368 : OAI22_X1 port map( A1 => n17177, A2 => n17285, B1 => n12828, B2 => 
                           n15141, ZN => n2265);
   U15369 : OAI22_X1 port map( A1 => n17178, A2 => n17288, B1 => n12827, B2 => 
                           n15141, ZN => n2266);
   U15370 : OAI22_X1 port map( A1 => n17178, A2 => n17300, B1 => n12826, B2 => 
                           n15141, ZN => n2267);
   U15371 : OAI22_X1 port map( A1 => n17140, A2 => n17270, B1 => n12961, B2 => 
                           n15148, ZN => n2132);
   U15372 : OAI22_X1 port map( A1 => n17141, A2 => n17273, B1 => n12960, B2 => 
                           n15148, ZN => n2133);
   U15373 : OAI22_X1 port map( A1 => n17141, A2 => n17276, B1 => n12959, B2 => 
                           n15148, ZN => n2134);
   U15374 : OAI22_X1 port map( A1 => n17141, A2 => n17279, B1 => n12958, B2 => 
                           n15148, ZN => n2135);
   U15375 : OAI22_X1 port map( A1 => n17141, A2 => n17282, B1 => n12957, B2 => 
                           n15148, ZN => n2136);
   U15376 : OAI22_X1 port map( A1 => n17141, A2 => n17285, B1 => n12956, B2 => 
                           n15148, ZN => n2137);
   U15377 : OAI22_X1 port map( A1 => n17142, A2 => n17288, B1 => n12955, B2 => 
                           n15148, ZN => n2138);
   U15378 : OAI22_X1 port map( A1 => n17142, A2 => n17300, B1 => n12954, B2 => 
                           n15148, ZN => n2139);
   U15379 : OAI22_X1 port map( A1 => n17104, A2 => n17270, B1 => n13089, B2 => 
                           n15153, ZN => n2004);
   U15380 : OAI22_X1 port map( A1 => n17105, A2 => n17273, B1 => n13088, B2 => 
                           n15153, ZN => n2005);
   U15381 : OAI22_X1 port map( A1 => n17105, A2 => n17276, B1 => n13087, B2 => 
                           n15153, ZN => n2006);
   U15382 : OAI22_X1 port map( A1 => n17105, A2 => n17279, B1 => n13086, B2 => 
                           n15153, ZN => n2007);
   U15383 : OAI22_X1 port map( A1 => n17105, A2 => n17282, B1 => n13085, B2 => 
                           n15153, ZN => n2008);
   U15384 : OAI22_X1 port map( A1 => n17105, A2 => n17285, B1 => n13084, B2 => 
                           n15153, ZN => n2009);
   U15385 : OAI22_X1 port map( A1 => n17106, A2 => n17288, B1 => n13083, B2 => 
                           n15153, ZN => n2010);
   U15386 : OAI22_X1 port map( A1 => n17106, A2 => n17300, B1 => n13082, B2 => 
                           n15153, ZN => n2011);
   U15387 : OAI22_X1 port map( A1 => n17068, A2 => n17271, B1 => n13217, B2 => 
                           n15158, ZN => n1876);
   U15388 : OAI22_X1 port map( A1 => n17069, A2 => n17274, B1 => n13216, B2 => 
                           n15158, ZN => n1877);
   U15389 : OAI22_X1 port map( A1 => n17069, A2 => n17277, B1 => n13215, B2 => 
                           n15158, ZN => n1878);
   U15390 : OAI22_X1 port map( A1 => n17069, A2 => n17280, B1 => n13214, B2 => 
                           n15158, ZN => n1879);
   U15391 : OAI22_X1 port map( A1 => n17069, A2 => n17283, B1 => n13213, B2 => 
                           n15158, ZN => n1880);
   U15392 : OAI22_X1 port map( A1 => n17069, A2 => n17286, B1 => n13212, B2 => 
                           n15158, ZN => n1881);
   U15393 : OAI22_X1 port map( A1 => n17070, A2 => n17289, B1 => n13211, B2 => 
                           n15158, ZN => n1882);
   U15394 : OAI22_X1 port map( A1 => n17070, A2 => n17301, B1 => n13210, B2 => 
                           n15158, ZN => n1883);
   U15395 : OAI22_X1 port map( A1 => n17059, A2 => n17271, B1 => n13249, B2 => 
                           n15159, ZN => n1844);
   U15396 : OAI22_X1 port map( A1 => n17060, A2 => n17274, B1 => n13248, B2 => 
                           n15159, ZN => n1845);
   U15397 : OAI22_X1 port map( A1 => n17060, A2 => n17277, B1 => n13247, B2 => 
                           n15159, ZN => n1846);
   U15398 : OAI22_X1 port map( A1 => n17060, A2 => n17280, B1 => n13246, B2 => 
                           n15159, ZN => n1847);
   U15399 : OAI22_X1 port map( A1 => n17060, A2 => n17283, B1 => n13245, B2 => 
                           n15159, ZN => n1848);
   U15400 : OAI22_X1 port map( A1 => n17060, A2 => n17286, B1 => n13244, B2 => 
                           n15159, ZN => n1849);
   U15401 : OAI22_X1 port map( A1 => n17061, A2 => n17289, B1 => n13243, B2 => 
                           n15159, ZN => n1850);
   U15402 : OAI22_X1 port map( A1 => n17061, A2 => n17301, B1 => n13242, B2 => 
                           n15159, ZN => n1851);
   U15403 : OAI22_X1 port map( A1 => n17050, A2 => n17271, B1 => n13281, B2 => 
                           n15161, ZN => n1812);
   U15404 : OAI22_X1 port map( A1 => n17051, A2 => n17274, B1 => n13280, B2 => 
                           n15161, ZN => n1813);
   U15405 : OAI22_X1 port map( A1 => n17051, A2 => n17277, B1 => n13279, B2 => 
                           n15161, ZN => n1814);
   U15406 : OAI22_X1 port map( A1 => n17051, A2 => n17280, B1 => n13278, B2 => 
                           n15161, ZN => n1815);
   U15407 : OAI22_X1 port map( A1 => n17051, A2 => n17283, B1 => n13277, B2 => 
                           n15161, ZN => n1816);
   U15408 : OAI22_X1 port map( A1 => n17051, A2 => n17286, B1 => n13276, B2 => 
                           n15161, ZN => n1817);
   U15409 : OAI22_X1 port map( A1 => n17052, A2 => n17289, B1 => n13275, B2 => 
                           n15161, ZN => n1818);
   U15410 : OAI22_X1 port map( A1 => n17052, A2 => n17301, B1 => n13274, B2 => 
                           n15161, ZN => n1819);
   U15411 : OAI22_X1 port map( A1 => n17041, A2 => n17271, B1 => n13313, B2 => 
                           n15162, ZN => n1780);
   U15412 : OAI22_X1 port map( A1 => n17042, A2 => n17274, B1 => n13312, B2 => 
                           n15162, ZN => n1781);
   U15413 : OAI22_X1 port map( A1 => n17042, A2 => n17277, B1 => n13311, B2 => 
                           n15162, ZN => n1782);
   U15414 : OAI22_X1 port map( A1 => n17042, A2 => n17280, B1 => n13310, B2 => 
                           n15162, ZN => n1783);
   U15415 : OAI22_X1 port map( A1 => n17042, A2 => n17283, B1 => n13309, B2 => 
                           n15162, ZN => n1784);
   U15416 : OAI22_X1 port map( A1 => n17042, A2 => n17286, B1 => n13308, B2 => 
                           n15162, ZN => n1785);
   U15417 : OAI22_X1 port map( A1 => n17043, A2 => n17289, B1 => n13307, B2 => 
                           n15162, ZN => n1786);
   U15418 : OAI22_X1 port map( A1 => n17043, A2 => n17301, B1 => n13306, B2 => 
                           n15162, ZN => n1787);
   U15419 : OAI22_X1 port map( A1 => n17032, A2 => n17271, B1 => n13345, B2 => 
                           n15163, ZN => n1748);
   U15420 : OAI22_X1 port map( A1 => n17033, A2 => n17274, B1 => n13344, B2 => 
                           n15163, ZN => n1749);
   U15421 : OAI22_X1 port map( A1 => n17033, A2 => n17277, B1 => n13343, B2 => 
                           n15163, ZN => n1750);
   U15422 : OAI22_X1 port map( A1 => n17033, A2 => n17280, B1 => n13342, B2 => 
                           n15163, ZN => n1751);
   U15423 : OAI22_X1 port map( A1 => n17033, A2 => n17283, B1 => n13341, B2 => 
                           n15163, ZN => n1752);
   U15424 : OAI22_X1 port map( A1 => n17033, A2 => n17286, B1 => n13340, B2 => 
                           n15163, ZN => n1753);
   U15425 : OAI22_X1 port map( A1 => n17034, A2 => n17289, B1 => n13339, B2 => 
                           n15163, ZN => n1754);
   U15426 : OAI22_X1 port map( A1 => n17034, A2 => n17301, B1 => n13338, B2 => 
                           n15163, ZN => n1755);
   U15427 : OAI22_X1 port map( A1 => n17023, A2 => n17271, B1 => n13377, B2 => 
                           n15165, ZN => n1716);
   U15428 : OAI22_X1 port map( A1 => n17024, A2 => n17274, B1 => n13376, B2 => 
                           n15165, ZN => n1717);
   U15429 : OAI22_X1 port map( A1 => n17024, A2 => n17277, B1 => n13375, B2 => 
                           n15165, ZN => n1718);
   U15430 : OAI22_X1 port map( A1 => n17024, A2 => n17280, B1 => n13374, B2 => 
                           n15165, ZN => n1719);
   U15431 : OAI22_X1 port map( A1 => n17024, A2 => n17283, B1 => n13373, B2 => 
                           n15165, ZN => n1720);
   U15432 : OAI22_X1 port map( A1 => n17024, A2 => n17286, B1 => n13372, B2 => 
                           n15165, ZN => n1721);
   U15433 : OAI22_X1 port map( A1 => n17025, A2 => n17289, B1 => n13371, B2 => 
                           n15165, ZN => n1722);
   U15434 : OAI22_X1 port map( A1 => n17025, A2 => n17301, B1 => n13370, B2 => 
                           n15165, ZN => n1723);
   U15435 : OAI22_X1 port map( A1 => n17014, A2 => n17271, B1 => n13409, B2 => 
                           n15167, ZN => n1684);
   U15436 : OAI22_X1 port map( A1 => n17015, A2 => n17274, B1 => n13408, B2 => 
                           n15167, ZN => n1685);
   U15437 : OAI22_X1 port map( A1 => n17015, A2 => n17277, B1 => n13407, B2 => 
                           n15167, ZN => n1686);
   U15438 : OAI22_X1 port map( A1 => n17015, A2 => n17280, B1 => n13406, B2 => 
                           n15167, ZN => n1687);
   U15439 : OAI22_X1 port map( A1 => n17015, A2 => n17283, B1 => n13405, B2 => 
                           n15167, ZN => n1688);
   U15440 : OAI22_X1 port map( A1 => n17015, A2 => n17286, B1 => n13404, B2 => 
                           n15167, ZN => n1689);
   U15441 : OAI22_X1 port map( A1 => n17016, A2 => n17289, B1 => n13403, B2 => 
                           n15167, ZN => n1690);
   U15442 : OAI22_X1 port map( A1 => n17016, A2 => n17301, B1 => n13402, B2 => 
                           n15167, ZN => n1691);
   U15443 : OAI22_X1 port map( A1 => n17005, A2 => n17271, B1 => n13441, B2 => 
                           n15168, ZN => n1652);
   U15444 : OAI22_X1 port map( A1 => n17006, A2 => n17274, B1 => n13440, B2 => 
                           n15168, ZN => n1653);
   U15445 : OAI22_X1 port map( A1 => n17006, A2 => n17277, B1 => n13439, B2 => 
                           n15168, ZN => n1654);
   U15446 : OAI22_X1 port map( A1 => n17006, A2 => n17280, B1 => n13438, B2 => 
                           n15168, ZN => n1655);
   U15447 : OAI22_X1 port map( A1 => n17006, A2 => n17283, B1 => n13437, B2 => 
                           n15168, ZN => n1656);
   U15448 : OAI22_X1 port map( A1 => n17006, A2 => n17286, B1 => n13436, B2 => 
                           n15168, ZN => n1657);
   U15449 : OAI22_X1 port map( A1 => n17007, A2 => n17289, B1 => n13435, B2 => 
                           n15168, ZN => n1658);
   U15450 : OAI22_X1 port map( A1 => n17007, A2 => n17301, B1 => n13434, B2 => 
                           n15168, ZN => n1659);
   U15451 : OAI22_X1 port map( A1 => n16996, A2 => n17271, B1 => n13473, B2 => 
                           n15169, ZN => n1620);
   U15452 : OAI22_X1 port map( A1 => n16997, A2 => n17274, B1 => n13472, B2 => 
                           n15169, ZN => n1621);
   U15453 : OAI22_X1 port map( A1 => n16997, A2 => n17277, B1 => n13471, B2 => 
                           n15169, ZN => n1622);
   U15454 : OAI22_X1 port map( A1 => n16997, A2 => n17280, B1 => n13470, B2 => 
                           n15169, ZN => n1623);
   U15455 : OAI22_X1 port map( A1 => n16997, A2 => n17283, B1 => n13469, B2 => 
                           n15169, ZN => n1624);
   U15456 : OAI22_X1 port map( A1 => n16997, A2 => n17286, B1 => n13468, B2 => 
                           n15169, ZN => n1625);
   U15457 : OAI22_X1 port map( A1 => n16998, A2 => n17289, B1 => n13467, B2 => 
                           n15169, ZN => n1626);
   U15458 : OAI22_X1 port map( A1 => n16998, A2 => n17301, B1 => n13466, B2 => 
                           n15169, ZN => n1627);
   U15459 : OAI22_X1 port map( A1 => n16987, A2 => n17272, B1 => n13505, B2 => 
                           n15170, ZN => n1588);
   U15460 : OAI22_X1 port map( A1 => n16988, A2 => n17275, B1 => n13504, B2 => 
                           n15170, ZN => n1589);
   U15461 : OAI22_X1 port map( A1 => n16988, A2 => n17278, B1 => n13503, B2 => 
                           n15170, ZN => n1590);
   U15462 : OAI22_X1 port map( A1 => n16988, A2 => n17281, B1 => n13502, B2 => 
                           n15170, ZN => n1591);
   U15463 : OAI22_X1 port map( A1 => n16988, A2 => n17284, B1 => n13501, B2 => 
                           n15170, ZN => n1592);
   U15464 : OAI22_X1 port map( A1 => n16988, A2 => n17287, B1 => n13500, B2 => 
                           n15170, ZN => n1593);
   U15465 : OAI22_X1 port map( A1 => n16989, A2 => n17290, B1 => n13499, B2 => 
                           n15170, ZN => n1594);
   U15466 : OAI22_X1 port map( A1 => n16989, A2 => n17302, B1 => n13498, B2 => 
                           n15170, ZN => n1595);
   U15467 : OAI22_X1 port map( A1 => n16978, A2 => n17272, B1 => n13537, B2 => 
                           n15172, ZN => n1556);
   U15468 : OAI22_X1 port map( A1 => n16979, A2 => n17275, B1 => n13536, B2 => 
                           n15172, ZN => n1557);
   U15469 : OAI22_X1 port map( A1 => n16979, A2 => n17278, B1 => n13535, B2 => 
                           n15172, ZN => n1558);
   U15470 : OAI22_X1 port map( A1 => n16979, A2 => n17281, B1 => n13534, B2 => 
                           n15172, ZN => n1559);
   U15471 : OAI22_X1 port map( A1 => n16979, A2 => n17284, B1 => n13533, B2 => 
                           n15172, ZN => n1560);
   U15472 : OAI22_X1 port map( A1 => n16979, A2 => n17287, B1 => n13532, B2 => 
                           n15172, ZN => n1561);
   U15473 : OAI22_X1 port map( A1 => n16980, A2 => n17290, B1 => n13531, B2 => 
                           n15172, ZN => n1562);
   U15474 : OAI22_X1 port map( A1 => n16980, A2 => n17302, B1 => n13530, B2 => 
                           n15172, ZN => n1563);
   U15475 : OAI22_X1 port map( A1 => n16969, A2 => n17272, B1 => n13569, B2 => 
                           n15173, ZN => n1524);
   U15476 : OAI22_X1 port map( A1 => n16970, A2 => n17275, B1 => n13568, B2 => 
                           n15173, ZN => n1525);
   U15477 : OAI22_X1 port map( A1 => n16970, A2 => n17278, B1 => n13567, B2 => 
                           n15173, ZN => n1526);
   U15478 : OAI22_X1 port map( A1 => n16970, A2 => n17281, B1 => n13566, B2 => 
                           n15173, ZN => n1527);
   U15479 : OAI22_X1 port map( A1 => n16970, A2 => n17284, B1 => n13565, B2 => 
                           n15173, ZN => n1528);
   U15480 : OAI22_X1 port map( A1 => n16970, A2 => n17287, B1 => n13564, B2 => 
                           n15173, ZN => n1529);
   U15481 : OAI22_X1 port map( A1 => n16971, A2 => n17290, B1 => n13563, B2 => 
                           n15173, ZN => n1530);
   U15482 : OAI22_X1 port map( A1 => n16971, A2 => n17302, B1 => n13562, B2 => 
                           n15173, ZN => n1531);
   U15483 : OAI22_X1 port map( A1 => n16960, A2 => n17272, B1 => n13601, B2 => 
                           n15174, ZN => n1492);
   U15484 : OAI22_X1 port map( A1 => n16961, A2 => n17275, B1 => n13600, B2 => 
                           n15174, ZN => n1493);
   U15485 : OAI22_X1 port map( A1 => n16961, A2 => n17278, B1 => n13599, B2 => 
                           n15174, ZN => n1494);
   U15486 : OAI22_X1 port map( A1 => n16961, A2 => n17281, B1 => n13598, B2 => 
                           n15174, ZN => n1495);
   U15487 : OAI22_X1 port map( A1 => n16961, A2 => n17284, B1 => n13597, B2 => 
                           n15174, ZN => n1496);
   U15488 : OAI22_X1 port map( A1 => n16961, A2 => n17287, B1 => n13596, B2 => 
                           n15174, ZN => n1497);
   U15489 : OAI22_X1 port map( A1 => n16962, A2 => n17290, B1 => n13595, B2 => 
                           n15174, ZN => n1498);
   U15490 : OAI22_X1 port map( A1 => n16962, A2 => n17302, B1 => n13594, B2 => 
                           n15174, ZN => n1499);
   U15491 : OAI22_X1 port map( A1 => n16951, A2 => n17272, B1 => n13633, B2 => 
                           n15175, ZN => n1460);
   U15492 : OAI22_X1 port map( A1 => n16952, A2 => n17275, B1 => n13632, B2 => 
                           n15175, ZN => n1461);
   U15493 : OAI22_X1 port map( A1 => n16952, A2 => n17278, B1 => n13631, B2 => 
                           n15175, ZN => n1462);
   U15494 : OAI22_X1 port map( A1 => n16952, A2 => n17281, B1 => n13630, B2 => 
                           n15175, ZN => n1463);
   U15495 : OAI22_X1 port map( A1 => n16952, A2 => n17284, B1 => n13629, B2 => 
                           n15175, ZN => n1464);
   U15496 : OAI22_X1 port map( A1 => n16952, A2 => n17287, B1 => n13628, B2 => 
                           n15175, ZN => n1465);
   U15497 : OAI22_X1 port map( A1 => n16953, A2 => n17290, B1 => n13627, B2 => 
                           n15175, ZN => n1466);
   U15498 : OAI22_X1 port map( A1 => n16953, A2 => n17302, B1 => n13626, B2 => 
                           n15175, ZN => n1467);
   U15499 : OAI22_X1 port map( A1 => n16942, A2 => n17272, B1 => n13665, B2 => 
                           n15177, ZN => n1428);
   U15500 : OAI22_X1 port map( A1 => n16943, A2 => n17275, B1 => n13664, B2 => 
                           n15177, ZN => n1429);
   U15501 : OAI22_X1 port map( A1 => n16943, A2 => n17278, B1 => n13663, B2 => 
                           n15177, ZN => n1430);
   U15502 : OAI22_X1 port map( A1 => n16943, A2 => n17281, B1 => n13662, B2 => 
                           n15177, ZN => n1431);
   U15503 : OAI22_X1 port map( A1 => n16943, A2 => n17284, B1 => n13661, B2 => 
                           n15177, ZN => n1432);
   U15504 : OAI22_X1 port map( A1 => n16943, A2 => n17287, B1 => n13660, B2 => 
                           n15177, ZN => n1433);
   U15505 : OAI22_X1 port map( A1 => n16944, A2 => n17290, B1 => n13659, B2 => 
                           n15177, ZN => n1434);
   U15506 : OAI22_X1 port map( A1 => n16944, A2 => n17302, B1 => n13658, B2 => 
                           n15177, ZN => n1435);
   U15507 : OAI22_X1 port map( A1 => n16933, A2 => n17272, B1 => n13697, B2 => 
                           n15178, ZN => n1396);
   U15508 : OAI22_X1 port map( A1 => n16934, A2 => n17275, B1 => n13696, B2 => 
                           n15178, ZN => n1397);
   U15509 : OAI22_X1 port map( A1 => n16934, A2 => n17278, B1 => n13695, B2 => 
                           n15178, ZN => n1398);
   U15510 : OAI22_X1 port map( A1 => n16934, A2 => n17281, B1 => n13694, B2 => 
                           n15178, ZN => n1399);
   U15511 : OAI22_X1 port map( A1 => n16934, A2 => n17284, B1 => n13693, B2 => 
                           n15178, ZN => n1400);
   U15512 : OAI22_X1 port map( A1 => n16934, A2 => n17287, B1 => n13692, B2 => 
                           n15178, ZN => n1401);
   U15513 : OAI22_X1 port map( A1 => n16935, A2 => n17290, B1 => n13691, B2 => 
                           n15178, ZN => n1402);
   U15514 : OAI22_X1 port map( A1 => n16935, A2 => n17302, B1 => n13690, B2 => 
                           n15178, ZN => n1403);
   U15515 : OAI221_X1 port map( B1 => n13528, B2 => n16774, C1 => n13592, C2 =>
                           n16771, A => n16314, ZN => n16312);
   U15516 : AOI22_X1 port map( A1 => n16768, A2 => n14979, B1 => n16767, B2 => 
                           n15003, ZN => n16314);
   U15517 : OAI221_X1 port map( B1 => n13527, B2 => n16774, C1 => n13591, C2 =>
                           n16771, A => n16297, ZN => n16295);
   U15518 : AOI22_X1 port map( A1 => n16768, A2 => n14978, B1 => n16767, B2 => 
                           n15002, ZN => n16297);
   U15519 : OAI221_X1 port map( B1 => n13526, B2 => n16774, C1 => n13590, C2 =>
                           n16771, A => n16280, ZN => n16278);
   U15520 : AOI22_X1 port map( A1 => n16768, A2 => n14977, B1 => n16767, B2 => 
                           n15001, ZN => n16280);
   U15521 : OAI221_X1 port map( B1 => n13525, B2 => n16774, C1 => n13589, C2 =>
                           n16771, A => n16263, ZN => n16261);
   U15522 : AOI22_X1 port map( A1 => n16768, A2 => n14976, B1 => n16767, B2 => 
                           n15000, ZN => n16263);
   U15523 : OAI221_X1 port map( B1 => n13524, B2 => n16774, C1 => n13588, C2 =>
                           n16771, A => n16246, ZN => n16244);
   U15524 : AOI22_X1 port map( A1 => n16768, A2 => n14975, B1 => n16767, B2 => 
                           n14999, ZN => n16246);
   U15525 : OAI221_X1 port map( B1 => n13523, B2 => n16774, C1 => n13587, C2 =>
                           n16771, A => n16229, ZN => n16227);
   U15526 : AOI22_X1 port map( A1 => n16768, A2 => n14974, B1 => n16767, B2 => 
                           n14998, ZN => n16229);
   U15527 : OAI221_X1 port map( B1 => n13522, B2 => n16774, C1 => n13586, C2 =>
                           n16771, A => n16212, ZN => n16210);
   U15528 : AOI22_X1 port map( A1 => n16768, A2 => n14973, B1 => n16767, B2 => 
                           n14997, ZN => n16212);
   U15529 : OAI221_X1 port map( B1 => n13521, B2 => n16774, C1 => n13585, C2 =>
                           n16771, A => n16195, ZN => n16193);
   U15530 : AOI22_X1 port map( A1 => n16768, A2 => n14972, B1 => n16766, B2 => 
                           n14996, ZN => n16195);
   U15531 : OAI221_X1 port map( B1 => n13505, B2 => n16776, C1 => n13569, C2 =>
                           n16773, A => n15923, ZN => n15921);
   U15532 : AOI22_X1 port map( A1 => n16770, A2 => n14868, B1 => n16765, B2 => 
                           n14876, ZN => n15923);
   U15533 : OAI221_X1 port map( B1 => n13697, B2 => n16797, C1 => n13409, C2 =>
                           n16794, A => n15920, ZN => n15916);
   U15534 : AOI22_X1 port map( A1 => n16791, A2 => n14852, B1 => n16786, B2 => 
                           n14860, ZN => n15920);
   U15535 : OAI221_X1 port map( B1 => n13504, B2 => n16776, C1 => n13568, C2 =>
                           n16773, A => n15906, ZN => n15904);
   U15536 : AOI22_X1 port map( A1 => n16770, A2 => n14867, B1 => n16765, B2 => 
                           n14875, ZN => n15906);
   U15537 : OAI221_X1 port map( B1 => n13696, B2 => n16797, C1 => n13408, C2 =>
                           n16794, A => n15903, ZN => n15899);
   U15538 : AOI22_X1 port map( A1 => n16791, A2 => n14851, B1 => n16786, B2 => 
                           n14859, ZN => n15903);
   U15539 : OAI221_X1 port map( B1 => n13503, B2 => n16776, C1 => n13567, C2 =>
                           n16773, A => n15889, ZN => n15887);
   U15540 : AOI22_X1 port map( A1 => n16770, A2 => n14866, B1 => n16765, B2 => 
                           n14874, ZN => n15889);
   U15541 : OAI221_X1 port map( B1 => n13695, B2 => n16797, C1 => n13407, C2 =>
                           n16794, A => n15886, ZN => n15882);
   U15542 : AOI22_X1 port map( A1 => n16791, A2 => n14850, B1 => n16786, B2 => 
                           n14858, ZN => n15886);
   U15543 : OAI221_X1 port map( B1 => n13502, B2 => n16776, C1 => n13566, C2 =>
                           n16773, A => n15872, ZN => n15870);
   U15544 : AOI22_X1 port map( A1 => n16770, A2 => n14865, B1 => n16765, B2 => 
                           n14873, ZN => n15872);
   U15545 : OAI221_X1 port map( B1 => n13694, B2 => n16797, C1 => n13406, C2 =>
                           n16794, A => n15869, ZN => n15865);
   U15546 : AOI22_X1 port map( A1 => n16791, A2 => n14849, B1 => n16786, B2 => 
                           n14857, ZN => n15869);
   U15547 : OAI221_X1 port map( B1 => n13501, B2 => n16776, C1 => n13565, C2 =>
                           n16773, A => n15855, ZN => n15853);
   U15548 : AOI22_X1 port map( A1 => n16770, A2 => n14864, B1 => n16765, B2 => 
                           n14872, ZN => n15855);
   U15549 : OAI221_X1 port map( B1 => n13693, B2 => n16797, C1 => n13405, C2 =>
                           n16794, A => n15852, ZN => n15848);
   U15550 : AOI22_X1 port map( A1 => n16791, A2 => n14848, B1 => n16786, B2 => 
                           n14856, ZN => n15852);
   U15551 : OAI221_X1 port map( B1 => n13500, B2 => n16776, C1 => n13564, C2 =>
                           n16773, A => n15838, ZN => n15836);
   U15552 : AOI22_X1 port map( A1 => n16770, A2 => n14863, B1 => n16765, B2 => 
                           n14871, ZN => n15838);
   U15553 : OAI221_X1 port map( B1 => n13692, B2 => n16797, C1 => n13404, C2 =>
                           n16794, A => n15835, ZN => n15831);
   U15554 : AOI22_X1 port map( A1 => n16791, A2 => n14847, B1 => n16786, B2 => 
                           n14855, ZN => n15835);
   U15555 : OAI221_X1 port map( B1 => n13499, B2 => n16776, C1 => n13563, C2 =>
                           n16773, A => n15821, ZN => n15819);
   U15556 : AOI22_X1 port map( A1 => n16770, A2 => n14862, B1 => n16765, B2 => 
                           n14870, ZN => n15821);
   U15557 : OAI221_X1 port map( B1 => n13691, B2 => n16797, C1 => n13403, C2 =>
                           n16794, A => n15818, ZN => n15814);
   U15558 : AOI22_X1 port map( A1 => n16791, A2 => n14846, B1 => n16786, B2 => 
                           n14854, ZN => n15818);
   U15559 : OAI221_X1 port map( B1 => n13498, B2 => n16776, C1 => n13562, C2 =>
                           n16773, A => n15790, ZN => n15784);
   U15560 : AOI22_X1 port map( A1 => n16770, A2 => n14861, B1 => n16765, B2 => 
                           n14869, ZN => n15790);
   U15561 : OAI221_X1 port map( B1 => n13690, B2 => n16797, C1 => n13402, C2 =>
                           n16794, A => n15780, ZN => n15765);
   U15562 : AOI22_X1 port map( A1 => n16791, A2 => n14845, B1 => n16786, B2 => 
                           n14853, ZN => n15780);
   U15563 : OAI221_X1 port map( B1 => n13528, B2 => n16867, C1 => n13592, C2 =>
                           n16864, A => n15733, ZN => n15731);
   U15564 : AOI22_X1 port map( A1 => n16861, A2 => n14979, B1 => n16860, B2 => 
                           n15003, ZN => n15733);
   U15565 : OAI221_X1 port map( B1 => n13527, B2 => n16867, C1 => n13591, C2 =>
                           n16864, A => n15716, ZN => n15714);
   U15566 : AOI22_X1 port map( A1 => n16861, A2 => n14978, B1 => n16860, B2 => 
                           n15002, ZN => n15716);
   U15567 : OAI221_X1 port map( B1 => n13526, B2 => n16867, C1 => n13590, C2 =>
                           n16864, A => n15699, ZN => n15697);
   U15568 : AOI22_X1 port map( A1 => n16861, A2 => n14977, B1 => n16860, B2 => 
                           n15001, ZN => n15699);
   U15569 : OAI221_X1 port map( B1 => n13525, B2 => n16867, C1 => n13589, C2 =>
                           n16864, A => n15682, ZN => n15680);
   U15570 : AOI22_X1 port map( A1 => n16861, A2 => n14976, B1 => n16860, B2 => 
                           n15000, ZN => n15682);
   U15571 : OAI221_X1 port map( B1 => n13524, B2 => n16867, C1 => n13588, C2 =>
                           n16864, A => n15665, ZN => n15663);
   U15572 : AOI22_X1 port map( A1 => n16861, A2 => n14975, B1 => n16860, B2 => 
                           n14999, ZN => n15665);
   U15573 : OAI221_X1 port map( B1 => n13523, B2 => n16867, C1 => n13587, C2 =>
                           n16864, A => n15648, ZN => n15646);
   U15574 : AOI22_X1 port map( A1 => n16861, A2 => n14974, B1 => n16860, B2 => 
                           n14998, ZN => n15648);
   U15575 : OAI221_X1 port map( B1 => n13522, B2 => n16867, C1 => n13586, C2 =>
                           n16864, A => n15631, ZN => n15629);
   U15576 : AOI22_X1 port map( A1 => n16861, A2 => n14973, B1 => n16860, B2 => 
                           n14997, ZN => n15631);
   U15577 : OAI221_X1 port map( B1 => n13521, B2 => n16867, C1 => n13585, C2 =>
                           n16864, A => n15614, ZN => n15612);
   U15578 : AOI22_X1 port map( A1 => n16861, A2 => n14972, B1 => n16859, B2 => 
                           n14996, ZN => n15614);
   U15579 : OAI221_X1 port map( B1 => n13505, B2 => n16869, C1 => n13569, C2 =>
                           n16866, A => n15342, ZN => n15340);
   U15580 : AOI22_X1 port map( A1 => n16863, A2 => n14868, B1 => n16858, B2 => 
                           n14876, ZN => n15342);
   U15581 : OAI221_X1 port map( B1 => n13697, B2 => n16890, C1 => n13409, C2 =>
                           n16887, A => n15339, ZN => n15335);
   U15582 : AOI22_X1 port map( A1 => n16884, A2 => n14852, B1 => n16879, B2 => 
                           n14860, ZN => n15339);
   U15583 : OAI221_X1 port map( B1 => n13504, B2 => n16869, C1 => n13568, C2 =>
                           n16866, A => n15325, ZN => n15323);
   U15584 : AOI22_X1 port map( A1 => n16863, A2 => n14867, B1 => n16858, B2 => 
                           n14875, ZN => n15325);
   U15585 : OAI221_X1 port map( B1 => n13696, B2 => n16890, C1 => n13408, C2 =>
                           n16887, A => n15322, ZN => n15318);
   U15586 : AOI22_X1 port map( A1 => n16884, A2 => n14851, B1 => n16879, B2 => 
                           n14859, ZN => n15322);
   U15587 : OAI221_X1 port map( B1 => n13503, B2 => n16869, C1 => n13567, C2 =>
                           n16866, A => n15308, ZN => n15306);
   U15588 : AOI22_X1 port map( A1 => n16863, A2 => n14866, B1 => n16858, B2 => 
                           n14874, ZN => n15308);
   U15589 : OAI221_X1 port map( B1 => n13695, B2 => n16890, C1 => n13407, C2 =>
                           n16887, A => n15305, ZN => n15301);
   U15590 : AOI22_X1 port map( A1 => n16884, A2 => n14850, B1 => n16879, B2 => 
                           n14858, ZN => n15305);
   U15591 : OAI221_X1 port map( B1 => n13502, B2 => n16869, C1 => n13566, C2 =>
                           n16866, A => n15291, ZN => n15289);
   U15592 : AOI22_X1 port map( A1 => n16863, A2 => n14865, B1 => n16858, B2 => 
                           n14873, ZN => n15291);
   U15593 : OAI221_X1 port map( B1 => n13694, B2 => n16890, C1 => n13406, C2 =>
                           n16887, A => n15288, ZN => n15284);
   U15594 : AOI22_X1 port map( A1 => n16884, A2 => n14849, B1 => n16879, B2 => 
                           n14857, ZN => n15288);
   U15595 : OAI221_X1 port map( B1 => n13501, B2 => n16869, C1 => n13565, C2 =>
                           n16866, A => n15274, ZN => n15272);
   U15596 : AOI22_X1 port map( A1 => n16863, A2 => n14864, B1 => n16858, B2 => 
                           n14872, ZN => n15274);
   U15597 : OAI221_X1 port map( B1 => n13693, B2 => n16890, C1 => n13405, C2 =>
                           n16887, A => n15271, ZN => n15267);
   U15598 : AOI22_X1 port map( A1 => n16884, A2 => n14848, B1 => n16879, B2 => 
                           n14856, ZN => n15271);
   U15599 : OAI221_X1 port map( B1 => n13500, B2 => n16869, C1 => n13564, C2 =>
                           n16866, A => n15257, ZN => n15255);
   U15600 : AOI22_X1 port map( A1 => n16863, A2 => n14863, B1 => n16858, B2 => 
                           n14871, ZN => n15257);
   U15601 : OAI221_X1 port map( B1 => n13692, B2 => n16890, C1 => n13404, C2 =>
                           n16887, A => n15254, ZN => n15250);
   U15602 : AOI22_X1 port map( A1 => n16884, A2 => n14847, B1 => n16879, B2 => 
                           n14855, ZN => n15254);
   U15603 : OAI221_X1 port map( B1 => n13499, B2 => n16869, C1 => n13563, C2 =>
                           n16866, A => n15240, ZN => n15238);
   U15604 : AOI22_X1 port map( A1 => n16863, A2 => n14862, B1 => n16858, B2 => 
                           n14870, ZN => n15240);
   U15605 : OAI221_X1 port map( B1 => n13691, B2 => n16890, C1 => n13403, C2 =>
                           n16887, A => n15237, ZN => n15233);
   U15606 : AOI22_X1 port map( A1 => n16884, A2 => n14846, B1 => n16879, B2 => 
                           n14854, ZN => n15237);
   U15607 : OAI221_X1 port map( B1 => n13498, B2 => n16869, C1 => n13562, C2 =>
                           n16866, A => n15209, ZN => n15203);
   U15608 : AOI22_X1 port map( A1 => n16863, A2 => n14861, B1 => n16858, B2 => 
                           n14869, ZN => n15209);
   U15609 : OAI221_X1 port map( B1 => n13690, B2 => n16890, C1 => n13402, C2 =>
                           n16887, A => n15199, ZN => n15184);
   U15610 : AOI22_X1 port map( A1 => n16884, A2 => n14845, B1 => n16879, B2 => 
                           n14853, ZN => n15199);
   U15611 : OAI22_X1 port map( A1 => n17127, A2 => n17198, B1 => n17126, B2 => 
                           n14685, ZN => n2076);
   U15612 : OAI22_X1 port map( A1 => n17127, A2 => n17201, B1 => n17126, B2 => 
                           n14684, ZN => n2077);
   U15613 : OAI22_X1 port map( A1 => n17127, A2 => n17204, B1 => n17126, B2 => 
                           n14683, ZN => n2078);
   U15614 : OAI22_X1 port map( A1 => n17127, A2 => n17207, B1 => n17126, B2 => 
                           n14682, ZN => n2079);
   U15615 : OAI22_X1 port map( A1 => n17127, A2 => n17210, B1 => n17126, B2 => 
                           n14681, ZN => n2080);
   U15616 : OAI22_X1 port map( A1 => n17128, A2 => n17213, B1 => n17126, B2 => 
                           n14680, ZN => n2081);
   U15617 : OAI22_X1 port map( A1 => n17128, A2 => n17216, B1 => n17126, B2 => 
                           n14679, ZN => n2082);
   U15618 : OAI22_X1 port map( A1 => n17128, A2 => n17219, B1 => n17126, B2 => 
                           n14678, ZN => n2083);
   U15619 : OAI22_X1 port map( A1 => n17128, A2 => n17222, B1 => n17126, B2 => 
                           n14677, ZN => n2084);
   U15620 : OAI22_X1 port map( A1 => n17128, A2 => n17225, B1 => n17126, B2 => 
                           n14676, ZN => n2085);
   U15621 : OAI22_X1 port map( A1 => n17129, A2 => n17228, B1 => n17126, B2 => 
                           n14675, ZN => n2086);
   U15622 : OAI22_X1 port map( A1 => n17129, A2 => n17231, B1 => n17126, B2 => 
                           n14674, ZN => n2087);
   U15623 : OAI22_X1 port map( A1 => n17129, A2 => n17234, B1 => n15149, B2 => 
                           n14673, ZN => n2088);
   U15624 : OAI22_X1 port map( A1 => n17129, A2 => n17237, B1 => n15149, B2 => 
                           n14672, ZN => n2089);
   U15625 : OAI22_X1 port map( A1 => n17129, A2 => n17240, B1 => n15149, B2 => 
                           n14671, ZN => n2090);
   U15626 : OAI22_X1 port map( A1 => n17130, A2 => n17243, B1 => n17126, B2 => 
                           n14670, ZN => n2091);
   U15627 : OAI22_X1 port map( A1 => n17130, A2 => n17246, B1 => n17126, B2 => 
                           n14669, ZN => n2092);
   U15628 : OAI22_X1 port map( A1 => n17130, A2 => n17249, B1 => n17126, B2 => 
                           n14668, ZN => n2093);
   U15629 : OAI22_X1 port map( A1 => n17130, A2 => n17252, B1 => n17126, B2 => 
                           n14667, ZN => n2094);
   U15630 : OAI22_X1 port map( A1 => n17130, A2 => n17255, B1 => n17126, B2 => 
                           n14666, ZN => n2095);
   U15631 : OAI22_X1 port map( A1 => n17131, A2 => n17258, B1 => n17126, B2 => 
                           n14665, ZN => n2096);
   U15632 : OAI22_X1 port map( A1 => n17131, A2 => n17261, B1 => n17126, B2 => 
                           n14664, ZN => n2097);
   U15633 : OAI22_X1 port map( A1 => n17131, A2 => n17264, B1 => n17126, B2 => 
                           n14663, ZN => n2098);
   U15634 : OAI22_X1 port map( A1 => n17131, A2 => n17267, B1 => n17126, B2 => 
                           n14662, ZN => n2099);
   U15635 : OAI22_X1 port map( A1 => n17181, A2 => n17198, B1 => n17180, B2 => 
                           n14557, ZN => n2268);
   U15636 : OAI22_X1 port map( A1 => n17181, A2 => n17201, B1 => n17180, B2 => 
                           n14556, ZN => n2269);
   U15637 : OAI22_X1 port map( A1 => n17181, A2 => n17204, B1 => n17180, B2 => 
                           n14555, ZN => n2270);
   U15638 : OAI22_X1 port map( A1 => n17181, A2 => n17207, B1 => n17180, B2 => 
                           n14554, ZN => n2271);
   U15639 : OAI22_X1 port map( A1 => n17181, A2 => n17210, B1 => n17180, B2 => 
                           n14553, ZN => n2272);
   U15640 : OAI22_X1 port map( A1 => n17182, A2 => n17213, B1 => n17180, B2 => 
                           n14552, ZN => n2273);
   U15641 : OAI22_X1 port map( A1 => n17182, A2 => n17216, B1 => n17180, B2 => 
                           n14551, ZN => n2274);
   U15642 : OAI22_X1 port map( A1 => n17182, A2 => n17219, B1 => n17180, B2 => 
                           n14550, ZN => n2275);
   U15643 : OAI22_X1 port map( A1 => n17182, A2 => n17222, B1 => n17180, B2 => 
                           n14549, ZN => n2276);
   U15644 : OAI22_X1 port map( A1 => n17182, A2 => n17225, B1 => n17180, B2 => 
                           n14548, ZN => n2277);
   U15645 : OAI22_X1 port map( A1 => n17183, A2 => n17228, B1 => n17180, B2 => 
                           n14547, ZN => n2278);
   U15646 : OAI22_X1 port map( A1 => n17183, A2 => n17231, B1 => n17180, B2 => 
                           n14546, ZN => n2279);
   U15647 : OAI22_X1 port map( A1 => n17183, A2 => n17234, B1 => n15139, B2 => 
                           n14545, ZN => n2280);
   U15648 : OAI22_X1 port map( A1 => n17183, A2 => n17237, B1 => n15139, B2 => 
                           n14544, ZN => n2281);
   U15649 : OAI22_X1 port map( A1 => n17183, A2 => n17240, B1 => n15139, B2 => 
                           n14543, ZN => n2282);
   U15650 : OAI22_X1 port map( A1 => n17184, A2 => n17243, B1 => n17180, B2 => 
                           n14542, ZN => n2283);
   U15651 : OAI22_X1 port map( A1 => n17184, A2 => n17246, B1 => n17180, B2 => 
                           n14541, ZN => n2284);
   U15652 : OAI22_X1 port map( A1 => n17184, A2 => n17249, B1 => n17180, B2 => 
                           n14540, ZN => n2285);
   U15653 : OAI22_X1 port map( A1 => n17184, A2 => n17252, B1 => n17180, B2 => 
                           n14539, ZN => n2286);
   U15654 : OAI22_X1 port map( A1 => n17184, A2 => n17255, B1 => n17180, B2 => 
                           n14538, ZN => n2287);
   U15655 : OAI22_X1 port map( A1 => n17185, A2 => n17258, B1 => n17180, B2 => 
                           n14537, ZN => n2288);
   U15656 : OAI22_X1 port map( A1 => n17185, A2 => n17261, B1 => n17180, B2 => 
                           n14536, ZN => n2289);
   U15657 : OAI22_X1 port map( A1 => n17185, A2 => n17264, B1 => n17180, B2 => 
                           n14535, ZN => n2290);
   U15658 : OAI22_X1 port map( A1 => n17185, A2 => n17267, B1 => n17180, B2 => 
                           n14534, ZN => n2291);
   U15659 : OAI22_X1 port map( A1 => n17190, A2 => n17198, B1 => n17189, B2 => 
                           n14525, ZN => n2300);
   U15660 : OAI22_X1 port map( A1 => n17190, A2 => n17201, B1 => n17189, B2 => 
                           n14524, ZN => n2301);
   U15661 : OAI22_X1 port map( A1 => n17190, A2 => n17204, B1 => n17189, B2 => 
                           n14523, ZN => n2302);
   U15662 : OAI22_X1 port map( A1 => n17190, A2 => n17207, B1 => n17189, B2 => 
                           n14522, ZN => n2303);
   U15663 : OAI22_X1 port map( A1 => n17190, A2 => n17210, B1 => n17189, B2 => 
                           n14521, ZN => n2304);
   U15664 : OAI22_X1 port map( A1 => n17191, A2 => n17213, B1 => n17189, B2 => 
                           n14520, ZN => n2305);
   U15665 : OAI22_X1 port map( A1 => n17191, A2 => n17216, B1 => n17189, B2 => 
                           n14519, ZN => n2306);
   U15666 : OAI22_X1 port map( A1 => n17191, A2 => n17219, B1 => n17189, B2 => 
                           n14518, ZN => n2307);
   U15667 : OAI22_X1 port map( A1 => n17191, A2 => n17222, B1 => n17189, B2 => 
                           n14517, ZN => n2308);
   U15668 : OAI22_X1 port map( A1 => n17191, A2 => n17225, B1 => n17189, B2 => 
                           n14516, ZN => n2309);
   U15669 : OAI22_X1 port map( A1 => n17192, A2 => n17228, B1 => n17189, B2 => 
                           n14515, ZN => n2310);
   U15670 : OAI22_X1 port map( A1 => n17192, A2 => n17231, B1 => n17189, B2 => 
                           n14514, ZN => n2311);
   U15671 : OAI22_X1 port map( A1 => n17192, A2 => n17234, B1 => n15137, B2 => 
                           n14513, ZN => n2312);
   U15672 : OAI22_X1 port map( A1 => n17192, A2 => n17237, B1 => n15137, B2 => 
                           n14512, ZN => n2313);
   U15673 : OAI22_X1 port map( A1 => n17192, A2 => n17240, B1 => n15137, B2 => 
                           n14511, ZN => n2314);
   U15674 : OAI22_X1 port map( A1 => n17193, A2 => n17243, B1 => n17189, B2 => 
                           n14510, ZN => n2315);
   U15675 : OAI22_X1 port map( A1 => n17193, A2 => n17246, B1 => n17189, B2 => 
                           n14509, ZN => n2316);
   U15676 : OAI22_X1 port map( A1 => n17193, A2 => n17249, B1 => n17189, B2 => 
                           n14508, ZN => n2317);
   U15677 : OAI22_X1 port map( A1 => n17193, A2 => n17252, B1 => n17189, B2 => 
                           n14507, ZN => n2318);
   U15678 : OAI22_X1 port map( A1 => n17193, A2 => n17255, B1 => n17189, B2 => 
                           n14506, ZN => n2319);
   U15679 : OAI22_X1 port map( A1 => n17194, A2 => n17258, B1 => n17189, B2 => 
                           n14505, ZN => n2320);
   U15680 : OAI22_X1 port map( A1 => n17194, A2 => n17261, B1 => n17189, B2 => 
                           n14504, ZN => n2321);
   U15681 : OAI22_X1 port map( A1 => n17194, A2 => n17264, B1 => n17189, B2 => 
                           n14503, ZN => n2322);
   U15682 : OAI22_X1 port map( A1 => n17194, A2 => n17267, B1 => n17189, B2 => 
                           n14502, ZN => n2323);
   U15683 : OAI22_X1 port map( A1 => n17292, A2 => n17198, B1 => n17291, B2 => 
                           n14493, ZN => n2332);
   U15684 : OAI22_X1 port map( A1 => n17292, A2 => n17201, B1 => n17291, B2 => 
                           n14492, ZN => n2333);
   U15685 : OAI22_X1 port map( A1 => n17292, A2 => n17204, B1 => n17291, B2 => 
                           n14491, ZN => n2334);
   U15686 : OAI22_X1 port map( A1 => n17292, A2 => n17207, B1 => n17291, B2 => 
                           n14490, ZN => n2335);
   U15687 : OAI22_X1 port map( A1 => n17292, A2 => n17210, B1 => n17291, B2 => 
                           n14489, ZN => n2336);
   U15688 : OAI22_X1 port map( A1 => n17293, A2 => n17213, B1 => n17291, B2 => 
                           n14488, ZN => n2337);
   U15689 : OAI22_X1 port map( A1 => n17293, A2 => n17216, B1 => n17291, B2 => 
                           n14487, ZN => n2338);
   U15690 : OAI22_X1 port map( A1 => n17293, A2 => n17219, B1 => n17291, B2 => 
                           n14486, ZN => n2339);
   U15691 : OAI22_X1 port map( A1 => n17293, A2 => n17222, B1 => n17291, B2 => 
                           n14485, ZN => n2340);
   U15692 : OAI22_X1 port map( A1 => n17293, A2 => n17225, B1 => n17291, B2 => 
                           n14484, ZN => n2341);
   U15693 : OAI22_X1 port map( A1 => n17294, A2 => n17228, B1 => n17291, B2 => 
                           n14483, ZN => n2342);
   U15694 : OAI22_X1 port map( A1 => n17294, A2 => n17231, B1 => n17291, B2 => 
                           n14482, ZN => n2343);
   U15695 : OAI22_X1 port map( A1 => n17294, A2 => n17234, B1 => n15103, B2 => 
                           n14481, ZN => n2344);
   U15696 : OAI22_X1 port map( A1 => n17294, A2 => n17237, B1 => n15103, B2 => 
                           n14480, ZN => n2345);
   U15697 : OAI22_X1 port map( A1 => n17294, A2 => n17240, B1 => n15103, B2 => 
                           n14479, ZN => n2346);
   U15698 : OAI22_X1 port map( A1 => n17295, A2 => n17243, B1 => n17291, B2 => 
                           n14478, ZN => n2347);
   U15699 : OAI22_X1 port map( A1 => n17295, A2 => n17246, B1 => n17291, B2 => 
                           n14477, ZN => n2348);
   U15700 : OAI22_X1 port map( A1 => n17295, A2 => n17249, B1 => n17291, B2 => 
                           n14476, ZN => n2349);
   U15701 : OAI22_X1 port map( A1 => n17295, A2 => n17252, B1 => n17291, B2 => 
                           n14475, ZN => n2350);
   U15702 : OAI22_X1 port map( A1 => n17295, A2 => n17255, B1 => n17291, B2 => 
                           n14474, ZN => n2351);
   U15703 : OAI22_X1 port map( A1 => n17296, A2 => n17258, B1 => n17291, B2 => 
                           n14473, ZN => n2352);
   U15704 : OAI22_X1 port map( A1 => n17296, A2 => n17261, B1 => n17291, B2 => 
                           n14472, ZN => n2353);
   U15705 : OAI22_X1 port map( A1 => n17296, A2 => n17264, B1 => n17291, B2 => 
                           n14471, ZN => n2354);
   U15706 : OAI22_X1 port map( A1 => n17296, A2 => n17267, B1 => n17291, B2 => 
                           n14470, ZN => n2355);
   U15707 : OAI22_X1 port map( A1 => n13753, A2 => n15179, B1 => n16919, B2 => 
                           n17200, ZN => n1340);
   U15708 : OAI22_X1 port map( A1 => n13752, A2 => n16918, B1 => n16919, B2 => 
                           n17203, ZN => n1341);
   U15709 : OAI22_X1 port map( A1 => n13751, A2 => n16918, B1 => n16919, B2 => 
                           n17206, ZN => n1342);
   U15710 : OAI22_X1 port map( A1 => n13750, A2 => n16918, B1 => n16919, B2 => 
                           n17209, ZN => n1343);
   U15711 : OAI22_X1 port map( A1 => n13749, A2 => n16918, B1 => n16920, B2 => 
                           n17212, ZN => n1344);
   U15712 : OAI22_X1 port map( A1 => n13748, A2 => n16918, B1 => n16920, B2 => 
                           n17215, ZN => n1345);
   U15713 : OAI22_X1 port map( A1 => n13747, A2 => n16918, B1 => n16920, B2 => 
                           n17218, ZN => n1346);
   U15714 : OAI22_X1 port map( A1 => n13746, A2 => n16918, B1 => n16920, B2 => 
                           n17221, ZN => n1347);
   U15715 : OAI22_X1 port map( A1 => n13745, A2 => n16918, B1 => n16921, B2 => 
                           n17224, ZN => n1348);
   U15716 : OAI22_X1 port map( A1 => n13744, A2 => n16918, B1 => n16921, B2 => 
                           n17227, ZN => n1349);
   U15717 : OAI22_X1 port map( A1 => n13743, A2 => n16918, B1 => n16921, B2 => 
                           n17230, ZN => n1350);
   U15718 : OAI22_X1 port map( A1 => n13742, A2 => n16918, B1 => n16921, B2 => 
                           n17233, ZN => n1351);
   U15719 : OAI22_X1 port map( A1 => n13741, A2 => n15179, B1 => n16922, B2 => 
                           n17236, ZN => n1352);
   U15720 : OAI22_X1 port map( A1 => n13740, A2 => n16918, B1 => n16922, B2 => 
                           n17239, ZN => n1353);
   U15721 : OAI22_X1 port map( A1 => n13739, A2 => n15179, B1 => n16922, B2 => 
                           n17242, ZN => n1354);
   U15722 : OAI22_X1 port map( A1 => n13738, A2 => n16918, B1 => n16922, B2 => 
                           n17245, ZN => n1355);
   U15723 : OAI22_X1 port map( A1 => n13737, A2 => n15179, B1 => n16923, B2 => 
                           n17248, ZN => n1356);
   U15724 : OAI22_X1 port map( A1 => n13736, A2 => n16918, B1 => n16923, B2 => 
                           n17251, ZN => n1357);
   U15725 : OAI22_X1 port map( A1 => n13735, A2 => n15179, B1 => n16923, B2 => 
                           n17254, ZN => n1358);
   U15726 : OAI22_X1 port map( A1 => n13734, A2 => n16918, B1 => n16923, B2 => 
                           n17257, ZN => n1359);
   U15727 : OAI22_X1 port map( A1 => n13733, A2 => n15179, B1 => n16924, B2 => 
                           n17260, ZN => n1360);
   U15728 : OAI22_X1 port map( A1 => n13732, A2 => n16918, B1 => n16924, B2 => 
                           n17263, ZN => n1361);
   U15729 : OAI22_X1 port map( A1 => n13731, A2 => n15179, B1 => n16924, B2 => 
                           n17266, ZN => n1362);
   U15730 : OAI22_X1 port map( A1 => n13730, A2 => n16918, B1 => n16924, B2 => 
                           n17269, ZN => n1363);
   U15731 : OAI22_X1 port map( A1 => n13729, A2 => n15179, B1 => n16925, B2 => 
                           n17272, ZN => n1364);
   U15732 : OAI22_X1 port map( A1 => n13728, A2 => n16918, B1 => n16925, B2 => 
                           n17275, ZN => n1365);
   U15733 : OAI22_X1 port map( A1 => n13727, A2 => n15179, B1 => n16925, B2 => 
                           n17278, ZN => n1366);
   U15734 : OAI22_X1 port map( A1 => n13726, A2 => n16918, B1 => n16925, B2 => 
                           n17281, ZN => n1367);
   U15735 : OAI22_X1 port map( A1 => n13725, A2 => n15179, B1 => n16926, B2 => 
                           n17284, ZN => n1368);
   U15736 : OAI22_X1 port map( A1 => n13724, A2 => n16918, B1 => n16926, B2 => 
                           n17287, ZN => n1369);
   U15737 : OAI22_X1 port map( A1 => n13723, A2 => n15179, B1 => n16926, B2 => 
                           n17290, ZN => n1370);
   U15738 : OAI22_X1 port map( A1 => n13722, A2 => n16918, B1 => n16926, B2 => 
                           n17302, ZN => n1371);
   U15739 : OAI22_X1 port map( A1 => n16983, A2 => n17200, B1 => n13529, B2 => 
                           n16982, ZN => n1564);
   U15740 : OAI22_X1 port map( A1 => n16983, A2 => n17203, B1 => n13528, B2 => 
                           n16982, ZN => n1565);
   U15741 : OAI22_X1 port map( A1 => n16983, A2 => n17206, B1 => n13527, B2 => 
                           n16982, ZN => n1566);
   U15742 : OAI22_X1 port map( A1 => n16983, A2 => n17209, B1 => n13526, B2 => 
                           n16982, ZN => n1567);
   U15743 : OAI22_X1 port map( A1 => n16983, A2 => n17212, B1 => n13525, B2 => 
                           n16982, ZN => n1568);
   U15744 : OAI22_X1 port map( A1 => n16984, A2 => n17215, B1 => n13524, B2 => 
                           n16982, ZN => n1569);
   U15745 : OAI22_X1 port map( A1 => n16984, A2 => n17218, B1 => n13523, B2 => 
                           n16982, ZN => n1570);
   U15746 : OAI22_X1 port map( A1 => n16984, A2 => n17221, B1 => n13522, B2 => 
                           n16982, ZN => n1571);
   U15747 : OAI22_X1 port map( A1 => n16984, A2 => n17224, B1 => n13521, B2 => 
                           n16982, ZN => n1572);
   U15748 : OAI22_X1 port map( A1 => n16984, A2 => n17227, B1 => n13520, B2 => 
                           n16982, ZN => n1573);
   U15749 : OAI22_X1 port map( A1 => n16985, A2 => n17230, B1 => n13519, B2 => 
                           n16982, ZN => n1574);
   U15750 : OAI22_X1 port map( A1 => n16985, A2 => n17233, B1 => n13518, B2 => 
                           n16982, ZN => n1575);
   U15751 : OAI22_X1 port map( A1 => n16985, A2 => n17236, B1 => n13517, B2 => 
                           n15170, ZN => n1576);
   U15752 : OAI22_X1 port map( A1 => n16985, A2 => n17239, B1 => n13516, B2 => 
                           n15170, ZN => n1577);
   U15753 : OAI22_X1 port map( A1 => n16985, A2 => n17242, B1 => n13515, B2 => 
                           n15170, ZN => n1578);
   U15754 : OAI22_X1 port map( A1 => n16986, A2 => n17245, B1 => n13514, B2 => 
                           n16982, ZN => n1579);
   U15755 : OAI22_X1 port map( A1 => n16986, A2 => n17248, B1 => n13513, B2 => 
                           n16982, ZN => n1580);
   U15756 : OAI22_X1 port map( A1 => n16986, A2 => n17251, B1 => n13512, B2 => 
                           n16982, ZN => n1581);
   U15757 : OAI22_X1 port map( A1 => n16986, A2 => n17254, B1 => n13511, B2 => 
                           n16982, ZN => n1582);
   U15758 : OAI22_X1 port map( A1 => n16986, A2 => n17257, B1 => n13510, B2 => 
                           n16982, ZN => n1583);
   U15759 : OAI22_X1 port map( A1 => n16987, A2 => n17260, B1 => n13509, B2 => 
                           n16982, ZN => n1584);
   U15760 : OAI22_X1 port map( A1 => n16987, A2 => n17263, B1 => n13508, B2 => 
                           n16982, ZN => n1585);
   U15761 : OAI22_X1 port map( A1 => n16987, A2 => n17266, B1 => n13507, B2 => 
                           n16982, ZN => n1586);
   U15762 : OAI22_X1 port map( A1 => n16987, A2 => n17269, B1 => n13506, B2 => 
                           n16982, ZN => n1587);
   U15763 : OAI22_X1 port map( A1 => n16929, A2 => n17200, B1 => n13721, B2 => 
                           n16928, ZN => n1372);
   U15764 : OAI22_X1 port map( A1 => n16929, A2 => n17203, B1 => n13720, B2 => 
                           n16928, ZN => n1373);
   U15765 : OAI22_X1 port map( A1 => n16929, A2 => n17206, B1 => n13719, B2 => 
                           n16928, ZN => n1374);
   U15766 : OAI22_X1 port map( A1 => n16929, A2 => n17209, B1 => n13718, B2 => 
                           n16928, ZN => n1375);
   U15767 : OAI22_X1 port map( A1 => n16929, A2 => n17212, B1 => n13717, B2 => 
                           n16928, ZN => n1376);
   U15768 : OAI22_X1 port map( A1 => n16930, A2 => n17215, B1 => n13716, B2 => 
                           n16928, ZN => n1377);
   U15769 : OAI22_X1 port map( A1 => n16930, A2 => n17218, B1 => n13715, B2 => 
                           n16928, ZN => n1378);
   U15770 : OAI22_X1 port map( A1 => n16930, A2 => n17221, B1 => n13714, B2 => 
                           n16928, ZN => n1379);
   U15771 : OAI22_X1 port map( A1 => n16930, A2 => n17224, B1 => n13713, B2 => 
                           n16928, ZN => n1380);
   U15772 : OAI22_X1 port map( A1 => n16930, A2 => n17227, B1 => n13712, B2 => 
                           n16928, ZN => n1381);
   U15773 : OAI22_X1 port map( A1 => n16931, A2 => n17230, B1 => n13711, B2 => 
                           n16928, ZN => n1382);
   U15774 : OAI22_X1 port map( A1 => n16931, A2 => n17233, B1 => n13710, B2 => 
                           n16928, ZN => n1383);
   U15775 : OAI22_X1 port map( A1 => n16931, A2 => n17236, B1 => n13709, B2 => 
                           n15178, ZN => n1384);
   U15776 : OAI22_X1 port map( A1 => n16931, A2 => n17239, B1 => n13708, B2 => 
                           n15178, ZN => n1385);
   U15777 : OAI22_X1 port map( A1 => n16931, A2 => n17242, B1 => n13707, B2 => 
                           n15178, ZN => n1386);
   U15778 : OAI22_X1 port map( A1 => n16932, A2 => n17245, B1 => n13706, B2 => 
                           n16928, ZN => n1387);
   U15779 : OAI22_X1 port map( A1 => n16932, A2 => n17248, B1 => n13705, B2 => 
                           n16928, ZN => n1388);
   U15780 : OAI22_X1 port map( A1 => n16932, A2 => n17251, B1 => n13704, B2 => 
                           n16928, ZN => n1389);
   U15781 : OAI22_X1 port map( A1 => n16932, A2 => n17254, B1 => n13703, B2 => 
                           n16928, ZN => n1390);
   U15782 : OAI22_X1 port map( A1 => n16932, A2 => n17257, B1 => n13702, B2 => 
                           n16928, ZN => n1391);
   U15783 : OAI22_X1 port map( A1 => n16933, A2 => n17260, B1 => n13701, B2 => 
                           n16928, ZN => n1392);
   U15784 : OAI22_X1 port map( A1 => n16933, A2 => n17263, B1 => n13700, B2 => 
                           n16928, ZN => n1393);
   U15785 : OAI22_X1 port map( A1 => n16933, A2 => n17266, B1 => n13699, B2 => 
                           n16928, ZN => n1394);
   U15786 : OAI22_X1 port map( A1 => n16933, A2 => n17269, B1 => n13698, B2 => 
                           n16928, ZN => n1395);
   U15787 : OAI22_X1 port map( A1 => n16974, A2 => n17200, B1 => n13561, B2 => 
                           n16973, ZN => n1532);
   U15788 : OAI22_X1 port map( A1 => n16974, A2 => n17203, B1 => n13560, B2 => 
                           n16973, ZN => n1533);
   U15789 : OAI22_X1 port map( A1 => n16974, A2 => n17206, B1 => n13559, B2 => 
                           n16973, ZN => n1534);
   U15790 : OAI22_X1 port map( A1 => n16974, A2 => n17209, B1 => n13558, B2 => 
                           n16973, ZN => n1535);
   U15791 : OAI22_X1 port map( A1 => n16974, A2 => n17212, B1 => n13557, B2 => 
                           n16973, ZN => n1536);
   U15792 : OAI22_X1 port map( A1 => n16975, A2 => n17215, B1 => n13556, B2 => 
                           n16973, ZN => n1537);
   U15793 : OAI22_X1 port map( A1 => n16975, A2 => n17218, B1 => n13555, B2 => 
                           n16973, ZN => n1538);
   U15794 : OAI22_X1 port map( A1 => n16975, A2 => n17221, B1 => n13554, B2 => 
                           n16973, ZN => n1539);
   U15795 : OAI22_X1 port map( A1 => n16975, A2 => n17224, B1 => n13553, B2 => 
                           n16973, ZN => n1540);
   U15796 : OAI22_X1 port map( A1 => n16975, A2 => n17227, B1 => n13552, B2 => 
                           n16973, ZN => n1541);
   U15797 : OAI22_X1 port map( A1 => n16976, A2 => n17230, B1 => n13551, B2 => 
                           n16973, ZN => n1542);
   U15798 : OAI22_X1 port map( A1 => n16976, A2 => n17233, B1 => n13550, B2 => 
                           n16973, ZN => n1543);
   U15799 : OAI22_X1 port map( A1 => n16976, A2 => n17236, B1 => n13549, B2 => 
                           n15172, ZN => n1544);
   U15800 : OAI22_X1 port map( A1 => n16976, A2 => n17239, B1 => n13548, B2 => 
                           n15172, ZN => n1545);
   U15801 : OAI22_X1 port map( A1 => n16976, A2 => n17242, B1 => n13547, B2 => 
                           n15172, ZN => n1546);
   U15802 : OAI22_X1 port map( A1 => n16977, A2 => n17245, B1 => n13546, B2 => 
                           n16973, ZN => n1547);
   U15803 : OAI22_X1 port map( A1 => n16977, A2 => n17248, B1 => n13545, B2 => 
                           n16973, ZN => n1548);
   U15804 : OAI22_X1 port map( A1 => n16977, A2 => n17251, B1 => n13544, B2 => 
                           n16973, ZN => n1549);
   U15805 : OAI22_X1 port map( A1 => n16977, A2 => n17254, B1 => n13543, B2 => 
                           n16973, ZN => n1550);
   U15806 : OAI22_X1 port map( A1 => n16977, A2 => n17257, B1 => n13542, B2 => 
                           n16973, ZN => n1551);
   U15807 : OAI22_X1 port map( A1 => n16978, A2 => n17260, B1 => n13541, B2 => 
                           n16973, ZN => n1552);
   U15808 : OAI22_X1 port map( A1 => n16978, A2 => n17263, B1 => n13540, B2 => 
                           n16973, ZN => n1553);
   U15809 : OAI22_X1 port map( A1 => n16978, A2 => n17266, B1 => n13539, B2 => 
                           n16973, ZN => n1554);
   U15810 : OAI22_X1 port map( A1 => n16978, A2 => n17269, B1 => n13538, B2 => 
                           n16973, ZN => n1555);
   U15811 : OAI22_X1 port map( A1 => n17172, A2 => n17198, B1 => n12857, B2 => 
                           n17171, ZN => n2236);
   U15812 : OAI22_X1 port map( A1 => n17172, A2 => n17201, B1 => n12856, B2 => 
                           n17171, ZN => n2237);
   U15813 : OAI22_X1 port map( A1 => n17172, A2 => n17204, B1 => n12855, B2 => 
                           n17171, ZN => n2238);
   U15814 : OAI22_X1 port map( A1 => n17172, A2 => n17207, B1 => n12854, B2 => 
                           n17171, ZN => n2239);
   U15815 : OAI22_X1 port map( A1 => n17172, A2 => n17210, B1 => n12853, B2 => 
                           n17171, ZN => n2240);
   U15816 : OAI22_X1 port map( A1 => n17173, A2 => n17213, B1 => n12852, B2 => 
                           n17171, ZN => n2241);
   U15817 : OAI22_X1 port map( A1 => n17173, A2 => n17216, B1 => n12851, B2 => 
                           n17171, ZN => n2242);
   U15818 : OAI22_X1 port map( A1 => n17173, A2 => n17219, B1 => n12850, B2 => 
                           n17171, ZN => n2243);
   U15819 : OAI22_X1 port map( A1 => n17173, A2 => n17222, B1 => n12849, B2 => 
                           n17171, ZN => n2244);
   U15820 : OAI22_X1 port map( A1 => n17173, A2 => n17225, B1 => n12848, B2 => 
                           n17171, ZN => n2245);
   U15821 : OAI22_X1 port map( A1 => n17174, A2 => n17228, B1 => n12847, B2 => 
                           n17171, ZN => n2246);
   U15822 : OAI22_X1 port map( A1 => n17174, A2 => n17231, B1 => n12846, B2 => 
                           n17171, ZN => n2247);
   U15823 : OAI22_X1 port map( A1 => n17174, A2 => n17234, B1 => n12845, B2 => 
                           n15141, ZN => n2248);
   U15824 : OAI22_X1 port map( A1 => n17174, A2 => n17237, B1 => n12844, B2 => 
                           n15141, ZN => n2249);
   U15825 : OAI22_X1 port map( A1 => n17174, A2 => n17240, B1 => n12843, B2 => 
                           n15141, ZN => n2250);
   U15826 : OAI22_X1 port map( A1 => n17175, A2 => n17243, B1 => n12842, B2 => 
                           n17171, ZN => n2251);
   U15827 : OAI22_X1 port map( A1 => n17175, A2 => n17246, B1 => n12841, B2 => 
                           n17171, ZN => n2252);
   U15828 : OAI22_X1 port map( A1 => n17175, A2 => n17249, B1 => n12840, B2 => 
                           n17171, ZN => n2253);
   U15829 : OAI22_X1 port map( A1 => n17175, A2 => n17252, B1 => n12839, B2 => 
                           n17171, ZN => n2254);
   U15830 : OAI22_X1 port map( A1 => n17175, A2 => n17255, B1 => n12838, B2 => 
                           n17171, ZN => n2255);
   U15831 : OAI22_X1 port map( A1 => n17176, A2 => n17258, B1 => n12837, B2 => 
                           n17171, ZN => n2256);
   U15832 : OAI22_X1 port map( A1 => n17176, A2 => n17261, B1 => n12836, B2 => 
                           n17171, ZN => n2257);
   U15833 : OAI22_X1 port map( A1 => n17176, A2 => n17264, B1 => n12835, B2 => 
                           n17171, ZN => n2258);
   U15834 : OAI22_X1 port map( A1 => n17176, A2 => n17267, B1 => n12834, B2 => 
                           n17171, ZN => n2259);
   U15835 : OAI22_X1 port map( A1 => n17136, A2 => n17198, B1 => n12985, B2 => 
                           n17135, ZN => n2108);
   U15836 : OAI22_X1 port map( A1 => n17136, A2 => n17201, B1 => n12984, B2 => 
                           n17135, ZN => n2109);
   U15837 : OAI22_X1 port map( A1 => n17136, A2 => n17204, B1 => n12983, B2 => 
                           n17135, ZN => n2110);
   U15838 : OAI22_X1 port map( A1 => n17136, A2 => n17207, B1 => n12982, B2 => 
                           n17135, ZN => n2111);
   U15839 : OAI22_X1 port map( A1 => n17136, A2 => n17210, B1 => n12981, B2 => 
                           n17135, ZN => n2112);
   U15840 : OAI22_X1 port map( A1 => n17137, A2 => n17213, B1 => n12980, B2 => 
                           n17135, ZN => n2113);
   U15841 : OAI22_X1 port map( A1 => n17137, A2 => n17216, B1 => n12979, B2 => 
                           n17135, ZN => n2114);
   U15842 : OAI22_X1 port map( A1 => n17137, A2 => n17219, B1 => n12978, B2 => 
                           n17135, ZN => n2115);
   U15843 : OAI22_X1 port map( A1 => n17137, A2 => n17222, B1 => n12977, B2 => 
                           n17135, ZN => n2116);
   U15844 : OAI22_X1 port map( A1 => n17137, A2 => n17225, B1 => n12976, B2 => 
                           n17135, ZN => n2117);
   U15845 : OAI22_X1 port map( A1 => n17138, A2 => n17228, B1 => n12975, B2 => 
                           n17135, ZN => n2118);
   U15846 : OAI22_X1 port map( A1 => n17138, A2 => n17231, B1 => n12974, B2 => 
                           n17135, ZN => n2119);
   U15847 : OAI22_X1 port map( A1 => n17138, A2 => n17234, B1 => n12973, B2 => 
                           n15148, ZN => n2120);
   U15848 : OAI22_X1 port map( A1 => n17138, A2 => n17237, B1 => n12972, B2 => 
                           n15148, ZN => n2121);
   U15849 : OAI22_X1 port map( A1 => n17138, A2 => n17240, B1 => n12971, B2 => 
                           n15148, ZN => n2122);
   U15850 : OAI22_X1 port map( A1 => n17139, A2 => n17243, B1 => n12970, B2 => 
                           n17135, ZN => n2123);
   U15851 : OAI22_X1 port map( A1 => n17139, A2 => n17246, B1 => n12969, B2 => 
                           n17135, ZN => n2124);
   U15852 : OAI22_X1 port map( A1 => n17139, A2 => n17249, B1 => n12968, B2 => 
                           n17135, ZN => n2125);
   U15853 : OAI22_X1 port map( A1 => n17139, A2 => n17252, B1 => n12967, B2 => 
                           n17135, ZN => n2126);
   U15854 : OAI22_X1 port map( A1 => n17139, A2 => n17255, B1 => n12966, B2 => 
                           n17135, ZN => n2127);
   U15855 : OAI22_X1 port map( A1 => n17140, A2 => n17258, B1 => n12965, B2 => 
                           n17135, ZN => n2128);
   U15856 : OAI22_X1 port map( A1 => n17140, A2 => n17261, B1 => n12964, B2 => 
                           n17135, ZN => n2129);
   U15857 : OAI22_X1 port map( A1 => n17140, A2 => n17264, B1 => n12963, B2 => 
                           n17135, ZN => n2130);
   U15858 : OAI22_X1 port map( A1 => n17140, A2 => n17267, B1 => n12962, B2 => 
                           n17135, ZN => n2131);
   U15859 : OAI22_X1 port map( A1 => n17100, A2 => n17198, B1 => n13113, B2 => 
                           n17099, ZN => n1980);
   U15860 : OAI22_X1 port map( A1 => n17100, A2 => n17201, B1 => n13112, B2 => 
                           n17099, ZN => n1981);
   U15861 : OAI22_X1 port map( A1 => n17100, A2 => n17204, B1 => n13111, B2 => 
                           n17099, ZN => n1982);
   U15862 : OAI22_X1 port map( A1 => n17100, A2 => n17207, B1 => n13110, B2 => 
                           n17099, ZN => n1983);
   U15863 : OAI22_X1 port map( A1 => n17100, A2 => n17210, B1 => n13109, B2 => 
                           n17099, ZN => n1984);
   U15864 : OAI22_X1 port map( A1 => n17101, A2 => n17213, B1 => n13108, B2 => 
                           n17099, ZN => n1985);
   U15865 : OAI22_X1 port map( A1 => n17101, A2 => n17216, B1 => n13107, B2 => 
                           n17099, ZN => n1986);
   U15866 : OAI22_X1 port map( A1 => n17101, A2 => n17219, B1 => n13106, B2 => 
                           n17099, ZN => n1987);
   U15867 : OAI22_X1 port map( A1 => n17101, A2 => n17222, B1 => n13105, B2 => 
                           n17099, ZN => n1988);
   U15868 : OAI22_X1 port map( A1 => n17101, A2 => n17225, B1 => n13104, B2 => 
                           n17099, ZN => n1989);
   U15869 : OAI22_X1 port map( A1 => n17102, A2 => n17228, B1 => n13103, B2 => 
                           n17099, ZN => n1990);
   U15870 : OAI22_X1 port map( A1 => n17102, A2 => n17231, B1 => n13102, B2 => 
                           n17099, ZN => n1991);
   U15871 : OAI22_X1 port map( A1 => n17102, A2 => n17234, B1 => n13101, B2 => 
                           n15153, ZN => n1992);
   U15872 : OAI22_X1 port map( A1 => n17102, A2 => n17237, B1 => n13100, B2 => 
                           n15153, ZN => n1993);
   U15873 : OAI22_X1 port map( A1 => n17102, A2 => n17240, B1 => n13099, B2 => 
                           n15153, ZN => n1994);
   U15874 : OAI22_X1 port map( A1 => n17103, A2 => n17243, B1 => n13098, B2 => 
                           n17099, ZN => n1995);
   U15875 : OAI22_X1 port map( A1 => n17103, A2 => n17246, B1 => n13097, B2 => 
                           n17099, ZN => n1996);
   U15876 : OAI22_X1 port map( A1 => n17103, A2 => n17249, B1 => n13096, B2 => 
                           n17099, ZN => n1997);
   U15877 : OAI22_X1 port map( A1 => n17103, A2 => n17252, B1 => n13095, B2 => 
                           n17099, ZN => n1998);
   U15878 : OAI22_X1 port map( A1 => n17103, A2 => n17255, B1 => n13094, B2 => 
                           n17099, ZN => n1999);
   U15879 : OAI22_X1 port map( A1 => n17104, A2 => n17258, B1 => n13093, B2 => 
                           n17099, ZN => n2000);
   U15880 : OAI22_X1 port map( A1 => n17104, A2 => n17261, B1 => n13092, B2 => 
                           n17099, ZN => n2001);
   U15881 : OAI22_X1 port map( A1 => n17104, A2 => n17264, B1 => n13091, B2 => 
                           n17099, ZN => n2002);
   U15882 : OAI22_X1 port map( A1 => n17104, A2 => n17267, B1 => n13090, B2 => 
                           n17099, ZN => n2003);
   U15883 : OAI22_X1 port map( A1 => n17064, A2 => n17199, B1 => n13241, B2 => 
                           n17063, ZN => n1852);
   U15884 : OAI22_X1 port map( A1 => n17064, A2 => n17202, B1 => n13240, B2 => 
                           n17063, ZN => n1853);
   U15885 : OAI22_X1 port map( A1 => n17064, A2 => n17205, B1 => n13239, B2 => 
                           n17063, ZN => n1854);
   U15886 : OAI22_X1 port map( A1 => n17064, A2 => n17208, B1 => n13238, B2 => 
                           n17063, ZN => n1855);
   U15887 : OAI22_X1 port map( A1 => n17064, A2 => n17211, B1 => n13237, B2 => 
                           n17063, ZN => n1856);
   U15888 : OAI22_X1 port map( A1 => n17065, A2 => n17214, B1 => n13236, B2 => 
                           n17063, ZN => n1857);
   U15889 : OAI22_X1 port map( A1 => n17065, A2 => n17217, B1 => n13235, B2 => 
                           n17063, ZN => n1858);
   U15890 : OAI22_X1 port map( A1 => n17065, A2 => n17220, B1 => n13234, B2 => 
                           n17063, ZN => n1859);
   U15891 : OAI22_X1 port map( A1 => n17065, A2 => n17223, B1 => n13233, B2 => 
                           n17063, ZN => n1860);
   U15892 : OAI22_X1 port map( A1 => n17065, A2 => n17226, B1 => n13232, B2 => 
                           n17063, ZN => n1861);
   U15893 : OAI22_X1 port map( A1 => n17066, A2 => n17229, B1 => n13231, B2 => 
                           n17063, ZN => n1862);
   U15894 : OAI22_X1 port map( A1 => n17066, A2 => n17232, B1 => n13230, B2 => 
                           n17063, ZN => n1863);
   U15895 : OAI22_X1 port map( A1 => n17066, A2 => n17235, B1 => n13229, B2 => 
                           n15158, ZN => n1864);
   U15896 : OAI22_X1 port map( A1 => n17066, A2 => n17238, B1 => n13228, B2 => 
                           n15158, ZN => n1865);
   U15897 : OAI22_X1 port map( A1 => n17066, A2 => n17241, B1 => n13227, B2 => 
                           n15158, ZN => n1866);
   U15898 : OAI22_X1 port map( A1 => n17067, A2 => n17244, B1 => n13226, B2 => 
                           n17063, ZN => n1867);
   U15899 : OAI22_X1 port map( A1 => n17067, A2 => n17247, B1 => n13225, B2 => 
                           n17063, ZN => n1868);
   U15900 : OAI22_X1 port map( A1 => n17067, A2 => n17250, B1 => n13224, B2 => 
                           n17063, ZN => n1869);
   U15901 : OAI22_X1 port map( A1 => n17067, A2 => n17253, B1 => n13223, B2 => 
                           n17063, ZN => n1870);
   U15902 : OAI22_X1 port map( A1 => n17067, A2 => n17256, B1 => n13222, B2 => 
                           n17063, ZN => n1871);
   U15903 : OAI22_X1 port map( A1 => n17068, A2 => n17259, B1 => n13221, B2 => 
                           n17063, ZN => n1872);
   U15904 : OAI22_X1 port map( A1 => n17068, A2 => n17262, B1 => n13220, B2 => 
                           n17063, ZN => n1873);
   U15905 : OAI22_X1 port map( A1 => n17068, A2 => n17265, B1 => n13219, B2 => 
                           n17063, ZN => n1874);
   U15906 : OAI22_X1 port map( A1 => n17068, A2 => n17268, B1 => n13218, B2 => 
                           n17063, ZN => n1875);
   U15907 : OAI22_X1 port map( A1 => n17055, A2 => n17199, B1 => n13273, B2 => 
                           n17054, ZN => n1820);
   U15908 : OAI22_X1 port map( A1 => n17055, A2 => n17202, B1 => n13272, B2 => 
                           n17054, ZN => n1821);
   U15909 : OAI22_X1 port map( A1 => n17055, A2 => n17205, B1 => n13271, B2 => 
                           n17054, ZN => n1822);
   U15910 : OAI22_X1 port map( A1 => n17055, A2 => n17208, B1 => n13270, B2 => 
                           n17054, ZN => n1823);
   U15911 : OAI22_X1 port map( A1 => n17055, A2 => n17211, B1 => n13269, B2 => 
                           n17054, ZN => n1824);
   U15912 : OAI22_X1 port map( A1 => n17056, A2 => n17214, B1 => n13268, B2 => 
                           n17054, ZN => n1825);
   U15913 : OAI22_X1 port map( A1 => n17056, A2 => n17217, B1 => n13267, B2 => 
                           n17054, ZN => n1826);
   U15914 : OAI22_X1 port map( A1 => n17056, A2 => n17220, B1 => n13266, B2 => 
                           n17054, ZN => n1827);
   U15915 : OAI22_X1 port map( A1 => n17056, A2 => n17223, B1 => n13265, B2 => 
                           n17054, ZN => n1828);
   U15916 : OAI22_X1 port map( A1 => n17056, A2 => n17226, B1 => n13264, B2 => 
                           n17054, ZN => n1829);
   U15917 : OAI22_X1 port map( A1 => n17057, A2 => n17229, B1 => n13263, B2 => 
                           n17054, ZN => n1830);
   U15918 : OAI22_X1 port map( A1 => n17057, A2 => n17232, B1 => n13262, B2 => 
                           n17054, ZN => n1831);
   U15919 : OAI22_X1 port map( A1 => n17057, A2 => n17235, B1 => n13261, B2 => 
                           n15159, ZN => n1832);
   U15920 : OAI22_X1 port map( A1 => n17057, A2 => n17238, B1 => n13260, B2 => 
                           n15159, ZN => n1833);
   U15921 : OAI22_X1 port map( A1 => n17057, A2 => n17241, B1 => n13259, B2 => 
                           n15159, ZN => n1834);
   U15922 : OAI22_X1 port map( A1 => n17058, A2 => n17244, B1 => n13258, B2 => 
                           n17054, ZN => n1835);
   U15923 : OAI22_X1 port map( A1 => n17058, A2 => n17247, B1 => n13257, B2 => 
                           n17054, ZN => n1836);
   U15924 : OAI22_X1 port map( A1 => n17058, A2 => n17250, B1 => n13256, B2 => 
                           n17054, ZN => n1837);
   U15925 : OAI22_X1 port map( A1 => n17058, A2 => n17253, B1 => n13255, B2 => 
                           n17054, ZN => n1838);
   U15926 : OAI22_X1 port map( A1 => n17058, A2 => n17256, B1 => n13254, B2 => 
                           n17054, ZN => n1839);
   U15927 : OAI22_X1 port map( A1 => n17059, A2 => n17259, B1 => n13253, B2 => 
                           n17054, ZN => n1840);
   U15928 : OAI22_X1 port map( A1 => n17059, A2 => n17262, B1 => n13252, B2 => 
                           n17054, ZN => n1841);
   U15929 : OAI22_X1 port map( A1 => n17059, A2 => n17265, B1 => n13251, B2 => 
                           n17054, ZN => n1842);
   U15930 : OAI22_X1 port map( A1 => n17059, A2 => n17268, B1 => n13250, B2 => 
                           n17054, ZN => n1843);
   U15931 : OAI22_X1 port map( A1 => n17046, A2 => n17199, B1 => n13305, B2 => 
                           n17045, ZN => n1788);
   U15932 : OAI22_X1 port map( A1 => n17046, A2 => n17202, B1 => n13304, B2 => 
                           n17045, ZN => n1789);
   U15933 : OAI22_X1 port map( A1 => n17046, A2 => n17205, B1 => n13303, B2 => 
                           n17045, ZN => n1790);
   U15934 : OAI22_X1 port map( A1 => n17046, A2 => n17208, B1 => n13302, B2 => 
                           n17045, ZN => n1791);
   U15935 : OAI22_X1 port map( A1 => n17046, A2 => n17211, B1 => n13301, B2 => 
                           n17045, ZN => n1792);
   U15936 : OAI22_X1 port map( A1 => n17047, A2 => n17214, B1 => n13300, B2 => 
                           n17045, ZN => n1793);
   U15937 : OAI22_X1 port map( A1 => n17047, A2 => n17217, B1 => n13299, B2 => 
                           n17045, ZN => n1794);
   U15938 : OAI22_X1 port map( A1 => n17047, A2 => n17220, B1 => n13298, B2 => 
                           n17045, ZN => n1795);
   U15939 : OAI22_X1 port map( A1 => n17047, A2 => n17223, B1 => n13297, B2 => 
                           n17045, ZN => n1796);
   U15940 : OAI22_X1 port map( A1 => n17047, A2 => n17226, B1 => n13296, B2 => 
                           n17045, ZN => n1797);
   U15941 : OAI22_X1 port map( A1 => n17048, A2 => n17229, B1 => n13295, B2 => 
                           n17045, ZN => n1798);
   U15942 : OAI22_X1 port map( A1 => n17048, A2 => n17232, B1 => n13294, B2 => 
                           n17045, ZN => n1799);
   U15943 : OAI22_X1 port map( A1 => n17048, A2 => n17235, B1 => n13293, B2 => 
                           n15161, ZN => n1800);
   U15944 : OAI22_X1 port map( A1 => n17048, A2 => n17238, B1 => n13292, B2 => 
                           n15161, ZN => n1801);
   U15945 : OAI22_X1 port map( A1 => n17048, A2 => n17241, B1 => n13291, B2 => 
                           n15161, ZN => n1802);
   U15946 : OAI22_X1 port map( A1 => n17049, A2 => n17244, B1 => n13290, B2 => 
                           n17045, ZN => n1803);
   U15947 : OAI22_X1 port map( A1 => n17049, A2 => n17247, B1 => n13289, B2 => 
                           n17045, ZN => n1804);
   U15948 : OAI22_X1 port map( A1 => n17049, A2 => n17250, B1 => n13288, B2 => 
                           n17045, ZN => n1805);
   U15949 : OAI22_X1 port map( A1 => n17049, A2 => n17253, B1 => n13287, B2 => 
                           n17045, ZN => n1806);
   U15950 : OAI22_X1 port map( A1 => n17049, A2 => n17256, B1 => n13286, B2 => 
                           n17045, ZN => n1807);
   U15951 : OAI22_X1 port map( A1 => n17050, A2 => n17259, B1 => n13285, B2 => 
                           n17045, ZN => n1808);
   U15952 : OAI22_X1 port map( A1 => n17050, A2 => n17262, B1 => n13284, B2 => 
                           n17045, ZN => n1809);
   U15953 : OAI22_X1 port map( A1 => n17050, A2 => n17265, B1 => n13283, B2 => 
                           n17045, ZN => n1810);
   U15954 : OAI22_X1 port map( A1 => n17050, A2 => n17268, B1 => n13282, B2 => 
                           n17045, ZN => n1811);
   U15955 : OAI22_X1 port map( A1 => n17037, A2 => n17199, B1 => n13337, B2 => 
                           n17036, ZN => n1756);
   U15956 : OAI22_X1 port map( A1 => n17037, A2 => n17202, B1 => n13336, B2 => 
                           n17036, ZN => n1757);
   U15957 : OAI22_X1 port map( A1 => n17037, A2 => n17205, B1 => n13335, B2 => 
                           n17036, ZN => n1758);
   U15958 : OAI22_X1 port map( A1 => n17037, A2 => n17208, B1 => n13334, B2 => 
                           n17036, ZN => n1759);
   U15959 : OAI22_X1 port map( A1 => n17037, A2 => n17211, B1 => n13333, B2 => 
                           n17036, ZN => n1760);
   U15960 : OAI22_X1 port map( A1 => n17038, A2 => n17214, B1 => n13332, B2 => 
                           n17036, ZN => n1761);
   U15961 : OAI22_X1 port map( A1 => n17038, A2 => n17217, B1 => n13331, B2 => 
                           n17036, ZN => n1762);
   U15962 : OAI22_X1 port map( A1 => n17038, A2 => n17220, B1 => n13330, B2 => 
                           n17036, ZN => n1763);
   U15963 : OAI22_X1 port map( A1 => n17038, A2 => n17223, B1 => n13329, B2 => 
                           n17036, ZN => n1764);
   U15964 : OAI22_X1 port map( A1 => n17038, A2 => n17226, B1 => n13328, B2 => 
                           n17036, ZN => n1765);
   U15965 : OAI22_X1 port map( A1 => n17039, A2 => n17229, B1 => n13327, B2 => 
                           n17036, ZN => n1766);
   U15966 : OAI22_X1 port map( A1 => n17039, A2 => n17232, B1 => n13326, B2 => 
                           n17036, ZN => n1767);
   U15967 : OAI22_X1 port map( A1 => n17039, A2 => n17235, B1 => n13325, B2 => 
                           n15162, ZN => n1768);
   U15968 : OAI22_X1 port map( A1 => n17039, A2 => n17238, B1 => n13324, B2 => 
                           n15162, ZN => n1769);
   U15969 : OAI22_X1 port map( A1 => n17039, A2 => n17241, B1 => n13323, B2 => 
                           n15162, ZN => n1770);
   U15970 : OAI22_X1 port map( A1 => n17040, A2 => n17244, B1 => n13322, B2 => 
                           n17036, ZN => n1771);
   U15971 : OAI22_X1 port map( A1 => n17040, A2 => n17247, B1 => n13321, B2 => 
                           n17036, ZN => n1772);
   U15972 : OAI22_X1 port map( A1 => n17040, A2 => n17250, B1 => n13320, B2 => 
                           n17036, ZN => n1773);
   U15973 : OAI22_X1 port map( A1 => n17040, A2 => n17253, B1 => n13319, B2 => 
                           n17036, ZN => n1774);
   U15974 : OAI22_X1 port map( A1 => n17040, A2 => n17256, B1 => n13318, B2 => 
                           n17036, ZN => n1775);
   U15975 : OAI22_X1 port map( A1 => n17041, A2 => n17259, B1 => n13317, B2 => 
                           n17036, ZN => n1776);
   U15976 : OAI22_X1 port map( A1 => n17041, A2 => n17262, B1 => n13316, B2 => 
                           n17036, ZN => n1777);
   U15977 : OAI22_X1 port map( A1 => n17041, A2 => n17265, B1 => n13315, B2 => 
                           n17036, ZN => n1778);
   U15978 : OAI22_X1 port map( A1 => n17041, A2 => n17268, B1 => n13314, B2 => 
                           n17036, ZN => n1779);
   U15979 : OAI22_X1 port map( A1 => n17028, A2 => n17199, B1 => n13369, B2 => 
                           n17027, ZN => n1724);
   U15980 : OAI22_X1 port map( A1 => n17028, A2 => n17202, B1 => n13368, B2 => 
                           n17027, ZN => n1725);
   U15981 : OAI22_X1 port map( A1 => n17028, A2 => n17205, B1 => n13367, B2 => 
                           n17027, ZN => n1726);
   U15982 : OAI22_X1 port map( A1 => n17028, A2 => n17208, B1 => n13366, B2 => 
                           n17027, ZN => n1727);
   U15983 : OAI22_X1 port map( A1 => n17028, A2 => n17211, B1 => n13365, B2 => 
                           n17027, ZN => n1728);
   U15984 : OAI22_X1 port map( A1 => n17029, A2 => n17214, B1 => n13364, B2 => 
                           n17027, ZN => n1729);
   U15985 : OAI22_X1 port map( A1 => n17029, A2 => n17217, B1 => n13363, B2 => 
                           n17027, ZN => n1730);
   U15986 : OAI22_X1 port map( A1 => n17029, A2 => n17220, B1 => n13362, B2 => 
                           n17027, ZN => n1731);
   U15987 : OAI22_X1 port map( A1 => n17029, A2 => n17223, B1 => n13361, B2 => 
                           n17027, ZN => n1732);
   U15988 : OAI22_X1 port map( A1 => n17029, A2 => n17226, B1 => n13360, B2 => 
                           n17027, ZN => n1733);
   U15989 : OAI22_X1 port map( A1 => n17030, A2 => n17229, B1 => n13359, B2 => 
                           n17027, ZN => n1734);
   U15990 : OAI22_X1 port map( A1 => n17030, A2 => n17232, B1 => n13358, B2 => 
                           n17027, ZN => n1735);
   U15991 : OAI22_X1 port map( A1 => n17030, A2 => n17235, B1 => n13357, B2 => 
                           n15163, ZN => n1736);
   U15992 : OAI22_X1 port map( A1 => n17030, A2 => n17238, B1 => n13356, B2 => 
                           n15163, ZN => n1737);
   U15993 : OAI22_X1 port map( A1 => n17030, A2 => n17241, B1 => n13355, B2 => 
                           n15163, ZN => n1738);
   U15994 : OAI22_X1 port map( A1 => n17031, A2 => n17244, B1 => n13354, B2 => 
                           n17027, ZN => n1739);
   U15995 : OAI22_X1 port map( A1 => n17031, A2 => n17247, B1 => n13353, B2 => 
                           n17027, ZN => n1740);
   U15996 : OAI22_X1 port map( A1 => n17031, A2 => n17250, B1 => n13352, B2 => 
                           n17027, ZN => n1741);
   U15997 : OAI22_X1 port map( A1 => n17031, A2 => n17253, B1 => n13351, B2 => 
                           n17027, ZN => n1742);
   U15998 : OAI22_X1 port map( A1 => n17031, A2 => n17256, B1 => n13350, B2 => 
                           n17027, ZN => n1743);
   U15999 : OAI22_X1 port map( A1 => n17032, A2 => n17259, B1 => n13349, B2 => 
                           n17027, ZN => n1744);
   U16000 : OAI22_X1 port map( A1 => n17032, A2 => n17262, B1 => n13348, B2 => 
                           n17027, ZN => n1745);
   U16001 : OAI22_X1 port map( A1 => n17032, A2 => n17265, B1 => n13347, B2 => 
                           n17027, ZN => n1746);
   U16002 : OAI22_X1 port map( A1 => n17032, A2 => n17268, B1 => n13346, B2 => 
                           n17027, ZN => n1747);
   U16003 : OAI22_X1 port map( A1 => n17019, A2 => n17199, B1 => n13401, B2 => 
                           n17018, ZN => n1692);
   U16004 : OAI22_X1 port map( A1 => n17019, A2 => n17202, B1 => n13400, B2 => 
                           n17018, ZN => n1693);
   U16005 : OAI22_X1 port map( A1 => n17019, A2 => n17205, B1 => n13399, B2 => 
                           n17018, ZN => n1694);
   U16006 : OAI22_X1 port map( A1 => n17019, A2 => n17208, B1 => n13398, B2 => 
                           n17018, ZN => n1695);
   U16007 : OAI22_X1 port map( A1 => n17019, A2 => n17211, B1 => n13397, B2 => 
                           n17018, ZN => n1696);
   U16008 : OAI22_X1 port map( A1 => n17020, A2 => n17214, B1 => n13396, B2 => 
                           n17018, ZN => n1697);
   U16009 : OAI22_X1 port map( A1 => n17020, A2 => n17217, B1 => n13395, B2 => 
                           n17018, ZN => n1698);
   U16010 : OAI22_X1 port map( A1 => n17020, A2 => n17220, B1 => n13394, B2 => 
                           n17018, ZN => n1699);
   U16011 : OAI22_X1 port map( A1 => n17020, A2 => n17223, B1 => n13393, B2 => 
                           n17018, ZN => n1700);
   U16012 : OAI22_X1 port map( A1 => n17020, A2 => n17226, B1 => n13392, B2 => 
                           n17018, ZN => n1701);
   U16013 : OAI22_X1 port map( A1 => n17021, A2 => n17229, B1 => n13391, B2 => 
                           n17018, ZN => n1702);
   U16014 : OAI22_X1 port map( A1 => n17021, A2 => n17232, B1 => n13390, B2 => 
                           n17018, ZN => n1703);
   U16015 : OAI22_X1 port map( A1 => n17021, A2 => n17235, B1 => n13389, B2 => 
                           n15165, ZN => n1704);
   U16016 : OAI22_X1 port map( A1 => n17021, A2 => n17238, B1 => n13388, B2 => 
                           n15165, ZN => n1705);
   U16017 : OAI22_X1 port map( A1 => n17021, A2 => n17241, B1 => n13387, B2 => 
                           n15165, ZN => n1706);
   U16018 : OAI22_X1 port map( A1 => n17022, A2 => n17244, B1 => n13386, B2 => 
                           n17018, ZN => n1707);
   U16019 : OAI22_X1 port map( A1 => n17022, A2 => n17247, B1 => n13385, B2 => 
                           n17018, ZN => n1708);
   U16020 : OAI22_X1 port map( A1 => n17022, A2 => n17250, B1 => n13384, B2 => 
                           n17018, ZN => n1709);
   U16021 : OAI22_X1 port map( A1 => n17022, A2 => n17253, B1 => n13383, B2 => 
                           n17018, ZN => n1710);
   U16022 : OAI22_X1 port map( A1 => n17022, A2 => n17256, B1 => n13382, B2 => 
                           n17018, ZN => n1711);
   U16023 : OAI22_X1 port map( A1 => n17023, A2 => n17259, B1 => n13381, B2 => 
                           n17018, ZN => n1712);
   U16024 : OAI22_X1 port map( A1 => n17023, A2 => n17262, B1 => n13380, B2 => 
                           n17018, ZN => n1713);
   U16025 : OAI22_X1 port map( A1 => n17023, A2 => n17265, B1 => n13379, B2 => 
                           n17018, ZN => n1714);
   U16026 : OAI22_X1 port map( A1 => n17023, A2 => n17268, B1 => n13378, B2 => 
                           n17018, ZN => n1715);
   U16027 : OAI22_X1 port map( A1 => n17010, A2 => n17199, B1 => n13433, B2 => 
                           n17009, ZN => n1660);
   U16028 : OAI22_X1 port map( A1 => n17010, A2 => n17202, B1 => n13432, B2 => 
                           n17009, ZN => n1661);
   U16029 : OAI22_X1 port map( A1 => n17010, A2 => n17205, B1 => n13431, B2 => 
                           n17009, ZN => n1662);
   U16030 : OAI22_X1 port map( A1 => n17010, A2 => n17208, B1 => n13430, B2 => 
                           n17009, ZN => n1663);
   U16031 : OAI22_X1 port map( A1 => n17010, A2 => n17211, B1 => n13429, B2 => 
                           n17009, ZN => n1664);
   U16032 : OAI22_X1 port map( A1 => n17011, A2 => n17214, B1 => n13428, B2 => 
                           n17009, ZN => n1665);
   U16033 : OAI22_X1 port map( A1 => n17011, A2 => n17217, B1 => n13427, B2 => 
                           n17009, ZN => n1666);
   U16034 : OAI22_X1 port map( A1 => n17011, A2 => n17220, B1 => n13426, B2 => 
                           n17009, ZN => n1667);
   U16035 : OAI22_X1 port map( A1 => n17011, A2 => n17223, B1 => n13425, B2 => 
                           n17009, ZN => n1668);
   U16036 : OAI22_X1 port map( A1 => n17011, A2 => n17226, B1 => n13424, B2 => 
                           n17009, ZN => n1669);
   U16037 : OAI22_X1 port map( A1 => n17012, A2 => n17229, B1 => n13423, B2 => 
                           n17009, ZN => n1670);
   U16038 : OAI22_X1 port map( A1 => n17012, A2 => n17232, B1 => n13422, B2 => 
                           n17009, ZN => n1671);
   U16039 : OAI22_X1 port map( A1 => n17012, A2 => n17235, B1 => n13421, B2 => 
                           n15167, ZN => n1672);
   U16040 : OAI22_X1 port map( A1 => n17012, A2 => n17238, B1 => n13420, B2 => 
                           n15167, ZN => n1673);
   U16041 : OAI22_X1 port map( A1 => n17012, A2 => n17241, B1 => n13419, B2 => 
                           n15167, ZN => n1674);
   U16042 : OAI22_X1 port map( A1 => n17013, A2 => n17244, B1 => n13418, B2 => 
                           n17009, ZN => n1675);
   U16043 : OAI22_X1 port map( A1 => n17013, A2 => n17247, B1 => n13417, B2 => 
                           n17009, ZN => n1676);
   U16044 : OAI22_X1 port map( A1 => n17013, A2 => n17250, B1 => n13416, B2 => 
                           n17009, ZN => n1677);
   U16045 : OAI22_X1 port map( A1 => n17013, A2 => n17253, B1 => n13415, B2 => 
                           n17009, ZN => n1678);
   U16046 : OAI22_X1 port map( A1 => n17013, A2 => n17256, B1 => n13414, B2 => 
                           n17009, ZN => n1679);
   U16047 : OAI22_X1 port map( A1 => n17014, A2 => n17259, B1 => n13413, B2 => 
                           n17009, ZN => n1680);
   U16048 : OAI22_X1 port map( A1 => n17014, A2 => n17262, B1 => n13412, B2 => 
                           n17009, ZN => n1681);
   U16049 : OAI22_X1 port map( A1 => n17014, A2 => n17265, B1 => n13411, B2 => 
                           n17009, ZN => n1682);
   U16050 : OAI22_X1 port map( A1 => n17014, A2 => n17268, B1 => n13410, B2 => 
                           n17009, ZN => n1683);
   U16051 : OAI22_X1 port map( A1 => n17001, A2 => n17199, B1 => n13465, B2 => 
                           n17000, ZN => n1628);
   U16052 : OAI22_X1 port map( A1 => n17001, A2 => n17202, B1 => n13464, B2 => 
                           n17000, ZN => n1629);
   U16053 : OAI22_X1 port map( A1 => n17001, A2 => n17205, B1 => n13463, B2 => 
                           n17000, ZN => n1630);
   U16054 : OAI22_X1 port map( A1 => n17001, A2 => n17208, B1 => n13462, B2 => 
                           n17000, ZN => n1631);
   U16055 : OAI22_X1 port map( A1 => n17001, A2 => n17211, B1 => n13461, B2 => 
                           n17000, ZN => n1632);
   U16056 : OAI22_X1 port map( A1 => n17002, A2 => n17214, B1 => n13460, B2 => 
                           n17000, ZN => n1633);
   U16057 : OAI22_X1 port map( A1 => n17002, A2 => n17217, B1 => n13459, B2 => 
                           n17000, ZN => n1634);
   U16058 : OAI22_X1 port map( A1 => n17002, A2 => n17220, B1 => n13458, B2 => 
                           n17000, ZN => n1635);
   U16059 : OAI22_X1 port map( A1 => n17002, A2 => n17223, B1 => n13457, B2 => 
                           n17000, ZN => n1636);
   U16060 : OAI22_X1 port map( A1 => n17002, A2 => n17226, B1 => n13456, B2 => 
                           n17000, ZN => n1637);
   U16061 : OAI22_X1 port map( A1 => n17003, A2 => n17229, B1 => n13455, B2 => 
                           n17000, ZN => n1638);
   U16062 : OAI22_X1 port map( A1 => n17003, A2 => n17232, B1 => n13454, B2 => 
                           n17000, ZN => n1639);
   U16063 : OAI22_X1 port map( A1 => n17003, A2 => n17235, B1 => n13453, B2 => 
                           n15168, ZN => n1640);
   U16064 : OAI22_X1 port map( A1 => n17003, A2 => n17238, B1 => n13452, B2 => 
                           n15168, ZN => n1641);
   U16065 : OAI22_X1 port map( A1 => n17003, A2 => n17241, B1 => n13451, B2 => 
                           n15168, ZN => n1642);
   U16066 : OAI22_X1 port map( A1 => n17004, A2 => n17244, B1 => n13450, B2 => 
                           n17000, ZN => n1643);
   U16067 : OAI22_X1 port map( A1 => n17004, A2 => n17247, B1 => n13449, B2 => 
                           n17000, ZN => n1644);
   U16068 : OAI22_X1 port map( A1 => n17004, A2 => n17250, B1 => n13448, B2 => 
                           n17000, ZN => n1645);
   U16069 : OAI22_X1 port map( A1 => n17004, A2 => n17253, B1 => n13447, B2 => 
                           n17000, ZN => n1646);
   U16070 : OAI22_X1 port map( A1 => n17004, A2 => n17256, B1 => n13446, B2 => 
                           n17000, ZN => n1647);
   U16071 : OAI22_X1 port map( A1 => n17005, A2 => n17259, B1 => n13445, B2 => 
                           n17000, ZN => n1648);
   U16072 : OAI22_X1 port map( A1 => n17005, A2 => n17262, B1 => n13444, B2 => 
                           n17000, ZN => n1649);
   U16073 : OAI22_X1 port map( A1 => n17005, A2 => n17265, B1 => n13443, B2 => 
                           n17000, ZN => n1650);
   U16074 : OAI22_X1 port map( A1 => n17005, A2 => n17268, B1 => n13442, B2 => 
                           n17000, ZN => n1651);
   U16075 : OAI22_X1 port map( A1 => n16992, A2 => n17199, B1 => n13497, B2 => 
                           n16991, ZN => n1596);
   U16076 : OAI22_X1 port map( A1 => n16992, A2 => n17202, B1 => n13496, B2 => 
                           n16991, ZN => n1597);
   U16077 : OAI22_X1 port map( A1 => n16992, A2 => n17205, B1 => n13495, B2 => 
                           n16991, ZN => n1598);
   U16078 : OAI22_X1 port map( A1 => n16992, A2 => n17208, B1 => n13494, B2 => 
                           n16991, ZN => n1599);
   U16079 : OAI22_X1 port map( A1 => n16992, A2 => n17211, B1 => n13493, B2 => 
                           n16991, ZN => n1600);
   U16080 : OAI22_X1 port map( A1 => n16993, A2 => n17214, B1 => n13492, B2 => 
                           n16991, ZN => n1601);
   U16081 : OAI22_X1 port map( A1 => n16993, A2 => n17217, B1 => n13491, B2 => 
                           n16991, ZN => n1602);
   U16082 : OAI22_X1 port map( A1 => n16993, A2 => n17220, B1 => n13490, B2 => 
                           n16991, ZN => n1603);
   U16083 : OAI22_X1 port map( A1 => n16993, A2 => n17223, B1 => n13489, B2 => 
                           n16991, ZN => n1604);
   U16084 : OAI22_X1 port map( A1 => n16993, A2 => n17226, B1 => n13488, B2 => 
                           n16991, ZN => n1605);
   U16085 : OAI22_X1 port map( A1 => n16994, A2 => n17229, B1 => n13487, B2 => 
                           n16991, ZN => n1606);
   U16086 : OAI22_X1 port map( A1 => n16994, A2 => n17232, B1 => n13486, B2 => 
                           n16991, ZN => n1607);
   U16087 : OAI22_X1 port map( A1 => n16994, A2 => n17235, B1 => n13485, B2 => 
                           n15169, ZN => n1608);
   U16088 : OAI22_X1 port map( A1 => n16994, A2 => n17238, B1 => n13484, B2 => 
                           n15169, ZN => n1609);
   U16089 : OAI22_X1 port map( A1 => n16994, A2 => n17241, B1 => n13483, B2 => 
                           n15169, ZN => n1610);
   U16090 : OAI22_X1 port map( A1 => n16995, A2 => n17244, B1 => n13482, B2 => 
                           n16991, ZN => n1611);
   U16091 : OAI22_X1 port map( A1 => n16995, A2 => n17247, B1 => n13481, B2 => 
                           n16991, ZN => n1612);
   U16092 : OAI22_X1 port map( A1 => n16995, A2 => n17250, B1 => n13480, B2 => 
                           n16991, ZN => n1613);
   U16093 : OAI22_X1 port map( A1 => n16995, A2 => n17253, B1 => n13479, B2 => 
                           n16991, ZN => n1614);
   U16094 : OAI22_X1 port map( A1 => n16995, A2 => n17256, B1 => n13478, B2 => 
                           n16991, ZN => n1615);
   U16095 : OAI22_X1 port map( A1 => n16996, A2 => n17259, B1 => n13477, B2 => 
                           n16991, ZN => n1616);
   U16096 : OAI22_X1 port map( A1 => n16996, A2 => n17262, B1 => n13476, B2 => 
                           n16991, ZN => n1617);
   U16097 : OAI22_X1 port map( A1 => n16996, A2 => n17265, B1 => n13475, B2 => 
                           n16991, ZN => n1618);
   U16098 : OAI22_X1 port map( A1 => n16996, A2 => n17268, B1 => n13474, B2 => 
                           n16991, ZN => n1619);
   U16099 : OAI22_X1 port map( A1 => n16965, A2 => n17200, B1 => n13593, B2 => 
                           n16964, ZN => n1500);
   U16100 : OAI22_X1 port map( A1 => n16965, A2 => n17203, B1 => n13592, B2 => 
                           n16964, ZN => n1501);
   U16101 : OAI22_X1 port map( A1 => n16965, A2 => n17206, B1 => n13591, B2 => 
                           n16964, ZN => n1502);
   U16102 : OAI22_X1 port map( A1 => n16965, A2 => n17209, B1 => n13590, B2 => 
                           n16964, ZN => n1503);
   U16103 : OAI22_X1 port map( A1 => n16965, A2 => n17212, B1 => n13589, B2 => 
                           n16964, ZN => n1504);
   U16104 : OAI22_X1 port map( A1 => n16966, A2 => n17215, B1 => n13588, B2 => 
                           n16964, ZN => n1505);
   U16105 : OAI22_X1 port map( A1 => n16966, A2 => n17218, B1 => n13587, B2 => 
                           n16964, ZN => n1506);
   U16106 : OAI22_X1 port map( A1 => n16966, A2 => n17221, B1 => n13586, B2 => 
                           n16964, ZN => n1507);
   U16107 : OAI22_X1 port map( A1 => n16966, A2 => n17224, B1 => n13585, B2 => 
                           n16964, ZN => n1508);
   U16108 : OAI22_X1 port map( A1 => n16966, A2 => n17227, B1 => n13584, B2 => 
                           n16964, ZN => n1509);
   U16109 : OAI22_X1 port map( A1 => n16967, A2 => n17230, B1 => n13583, B2 => 
                           n16964, ZN => n1510);
   U16110 : OAI22_X1 port map( A1 => n16967, A2 => n17233, B1 => n13582, B2 => 
                           n16964, ZN => n1511);
   U16111 : OAI22_X1 port map( A1 => n16967, A2 => n17236, B1 => n13581, B2 => 
                           n15173, ZN => n1512);
   U16112 : OAI22_X1 port map( A1 => n16967, A2 => n17239, B1 => n13580, B2 => 
                           n15173, ZN => n1513);
   U16113 : OAI22_X1 port map( A1 => n16967, A2 => n17242, B1 => n13579, B2 => 
                           n15173, ZN => n1514);
   U16114 : OAI22_X1 port map( A1 => n16968, A2 => n17245, B1 => n13578, B2 => 
                           n16964, ZN => n1515);
   U16115 : OAI22_X1 port map( A1 => n16968, A2 => n17248, B1 => n13577, B2 => 
                           n16964, ZN => n1516);
   U16116 : OAI22_X1 port map( A1 => n16968, A2 => n17251, B1 => n13576, B2 => 
                           n16964, ZN => n1517);
   U16117 : OAI22_X1 port map( A1 => n16968, A2 => n17254, B1 => n13575, B2 => 
                           n16964, ZN => n1518);
   U16118 : OAI22_X1 port map( A1 => n16968, A2 => n17257, B1 => n13574, B2 => 
                           n16964, ZN => n1519);
   U16119 : OAI22_X1 port map( A1 => n16969, A2 => n17260, B1 => n13573, B2 => 
                           n16964, ZN => n1520);
   U16120 : OAI22_X1 port map( A1 => n16969, A2 => n17263, B1 => n13572, B2 => 
                           n16964, ZN => n1521);
   U16121 : OAI22_X1 port map( A1 => n16969, A2 => n17266, B1 => n13571, B2 => 
                           n16964, ZN => n1522);
   U16122 : OAI22_X1 port map( A1 => n16969, A2 => n17269, B1 => n13570, B2 => 
                           n16964, ZN => n1523);
   U16123 : OAI22_X1 port map( A1 => n16956, A2 => n17200, B1 => n13625, B2 => 
                           n16955, ZN => n1468);
   U16124 : OAI22_X1 port map( A1 => n16956, A2 => n17203, B1 => n13624, B2 => 
                           n16955, ZN => n1469);
   U16125 : OAI22_X1 port map( A1 => n16956, A2 => n17206, B1 => n13623, B2 => 
                           n16955, ZN => n1470);
   U16126 : OAI22_X1 port map( A1 => n16956, A2 => n17209, B1 => n13622, B2 => 
                           n16955, ZN => n1471);
   U16127 : OAI22_X1 port map( A1 => n16956, A2 => n17212, B1 => n13621, B2 => 
                           n16955, ZN => n1472);
   U16128 : OAI22_X1 port map( A1 => n16957, A2 => n17215, B1 => n13620, B2 => 
                           n16955, ZN => n1473);
   U16129 : OAI22_X1 port map( A1 => n16957, A2 => n17218, B1 => n13619, B2 => 
                           n16955, ZN => n1474);
   U16130 : OAI22_X1 port map( A1 => n16957, A2 => n17221, B1 => n13618, B2 => 
                           n16955, ZN => n1475);
   U16131 : OAI22_X1 port map( A1 => n16957, A2 => n17224, B1 => n13617, B2 => 
                           n16955, ZN => n1476);
   U16132 : OAI22_X1 port map( A1 => n16957, A2 => n17227, B1 => n13616, B2 => 
                           n16955, ZN => n1477);
   U16133 : OAI22_X1 port map( A1 => n16958, A2 => n17230, B1 => n13615, B2 => 
                           n16955, ZN => n1478);
   U16134 : OAI22_X1 port map( A1 => n16958, A2 => n17233, B1 => n13614, B2 => 
                           n16955, ZN => n1479);
   U16135 : OAI22_X1 port map( A1 => n16958, A2 => n17236, B1 => n13613, B2 => 
                           n15174, ZN => n1480);
   U16136 : OAI22_X1 port map( A1 => n16958, A2 => n17239, B1 => n13612, B2 => 
                           n15174, ZN => n1481);
   U16137 : OAI22_X1 port map( A1 => n16958, A2 => n17242, B1 => n13611, B2 => 
                           n15174, ZN => n1482);
   U16138 : OAI22_X1 port map( A1 => n16959, A2 => n17245, B1 => n13610, B2 => 
                           n16955, ZN => n1483);
   U16139 : OAI22_X1 port map( A1 => n16959, A2 => n17248, B1 => n13609, B2 => 
                           n16955, ZN => n1484);
   U16140 : OAI22_X1 port map( A1 => n16959, A2 => n17251, B1 => n13608, B2 => 
                           n16955, ZN => n1485);
   U16141 : OAI22_X1 port map( A1 => n16959, A2 => n17254, B1 => n13607, B2 => 
                           n16955, ZN => n1486);
   U16142 : OAI22_X1 port map( A1 => n16959, A2 => n17257, B1 => n13606, B2 => 
                           n16955, ZN => n1487);
   U16143 : OAI22_X1 port map( A1 => n16960, A2 => n17260, B1 => n13605, B2 => 
                           n16955, ZN => n1488);
   U16144 : OAI22_X1 port map( A1 => n16960, A2 => n17263, B1 => n13604, B2 => 
                           n16955, ZN => n1489);
   U16145 : OAI22_X1 port map( A1 => n16960, A2 => n17266, B1 => n13603, B2 => 
                           n16955, ZN => n1490);
   U16146 : OAI22_X1 port map( A1 => n16960, A2 => n17269, B1 => n13602, B2 => 
                           n16955, ZN => n1491);
   U16147 : OAI22_X1 port map( A1 => n16947, A2 => n17200, B1 => n13657, B2 => 
                           n16946, ZN => n1436);
   U16148 : OAI22_X1 port map( A1 => n16947, A2 => n17203, B1 => n13656, B2 => 
                           n16946, ZN => n1437);
   U16149 : OAI22_X1 port map( A1 => n16947, A2 => n17206, B1 => n13655, B2 => 
                           n16946, ZN => n1438);
   U16150 : OAI22_X1 port map( A1 => n16947, A2 => n17209, B1 => n13654, B2 => 
                           n16946, ZN => n1439);
   U16151 : OAI22_X1 port map( A1 => n16947, A2 => n17212, B1 => n13653, B2 => 
                           n16946, ZN => n1440);
   U16152 : OAI22_X1 port map( A1 => n16948, A2 => n17215, B1 => n13652, B2 => 
                           n16946, ZN => n1441);
   U16153 : OAI22_X1 port map( A1 => n16948, A2 => n17218, B1 => n13651, B2 => 
                           n16946, ZN => n1442);
   U16154 : OAI22_X1 port map( A1 => n16948, A2 => n17221, B1 => n13650, B2 => 
                           n16946, ZN => n1443);
   U16155 : OAI22_X1 port map( A1 => n16948, A2 => n17224, B1 => n13649, B2 => 
                           n16946, ZN => n1444);
   U16156 : OAI22_X1 port map( A1 => n16948, A2 => n17227, B1 => n13648, B2 => 
                           n16946, ZN => n1445);
   U16157 : OAI22_X1 port map( A1 => n16949, A2 => n17230, B1 => n13647, B2 => 
                           n16946, ZN => n1446);
   U16158 : OAI22_X1 port map( A1 => n16949, A2 => n17233, B1 => n13646, B2 => 
                           n16946, ZN => n1447);
   U16159 : OAI22_X1 port map( A1 => n16949, A2 => n17236, B1 => n13645, B2 => 
                           n15175, ZN => n1448);
   U16160 : OAI22_X1 port map( A1 => n16949, A2 => n17239, B1 => n13644, B2 => 
                           n15175, ZN => n1449);
   U16161 : OAI22_X1 port map( A1 => n16949, A2 => n17242, B1 => n13643, B2 => 
                           n15175, ZN => n1450);
   U16162 : OAI22_X1 port map( A1 => n16950, A2 => n17245, B1 => n13642, B2 => 
                           n16946, ZN => n1451);
   U16163 : OAI22_X1 port map( A1 => n16950, A2 => n17248, B1 => n13641, B2 => 
                           n16946, ZN => n1452);
   U16164 : OAI22_X1 port map( A1 => n16950, A2 => n17251, B1 => n13640, B2 => 
                           n16946, ZN => n1453);
   U16165 : OAI22_X1 port map( A1 => n16950, A2 => n17254, B1 => n13639, B2 => 
                           n16946, ZN => n1454);
   U16166 : OAI22_X1 port map( A1 => n16950, A2 => n17257, B1 => n13638, B2 => 
                           n16946, ZN => n1455);
   U16167 : OAI22_X1 port map( A1 => n16951, A2 => n17260, B1 => n13637, B2 => 
                           n16946, ZN => n1456);
   U16168 : OAI22_X1 port map( A1 => n16951, A2 => n17263, B1 => n13636, B2 => 
                           n16946, ZN => n1457);
   U16169 : OAI22_X1 port map( A1 => n16951, A2 => n17266, B1 => n13635, B2 => 
                           n16946, ZN => n1458);
   U16170 : OAI22_X1 port map( A1 => n16951, A2 => n17269, B1 => n13634, B2 => 
                           n16946, ZN => n1459);
   U16171 : OAI22_X1 port map( A1 => n16938, A2 => n17200, B1 => n13689, B2 => 
                           n16937, ZN => n1404);
   U16172 : OAI22_X1 port map( A1 => n16938, A2 => n17203, B1 => n13688, B2 => 
                           n16937, ZN => n1405);
   U16173 : OAI22_X1 port map( A1 => n16938, A2 => n17206, B1 => n13687, B2 => 
                           n16937, ZN => n1406);
   U16174 : OAI22_X1 port map( A1 => n16938, A2 => n17209, B1 => n13686, B2 => 
                           n16937, ZN => n1407);
   U16175 : OAI22_X1 port map( A1 => n16938, A2 => n17212, B1 => n13685, B2 => 
                           n16937, ZN => n1408);
   U16176 : OAI22_X1 port map( A1 => n16939, A2 => n17215, B1 => n13684, B2 => 
                           n16937, ZN => n1409);
   U16177 : OAI22_X1 port map( A1 => n16939, A2 => n17218, B1 => n13683, B2 => 
                           n16937, ZN => n1410);
   U16178 : OAI22_X1 port map( A1 => n16939, A2 => n17221, B1 => n13682, B2 => 
                           n16937, ZN => n1411);
   U16179 : OAI22_X1 port map( A1 => n16939, A2 => n17224, B1 => n13681, B2 => 
                           n16937, ZN => n1412);
   U16180 : OAI22_X1 port map( A1 => n16939, A2 => n17227, B1 => n13680, B2 => 
                           n16937, ZN => n1413);
   U16181 : OAI22_X1 port map( A1 => n16940, A2 => n17230, B1 => n13679, B2 => 
                           n16937, ZN => n1414);
   U16182 : OAI22_X1 port map( A1 => n16940, A2 => n17233, B1 => n13678, B2 => 
                           n16937, ZN => n1415);
   U16183 : OAI22_X1 port map( A1 => n16940, A2 => n17236, B1 => n13677, B2 => 
                           n15177, ZN => n1416);
   U16184 : OAI22_X1 port map( A1 => n16940, A2 => n17239, B1 => n13676, B2 => 
                           n15177, ZN => n1417);
   U16185 : OAI22_X1 port map( A1 => n16940, A2 => n17242, B1 => n13675, B2 => 
                           n15177, ZN => n1418);
   U16186 : OAI22_X1 port map( A1 => n16941, A2 => n17245, B1 => n13674, B2 => 
                           n16937, ZN => n1419);
   U16187 : OAI22_X1 port map( A1 => n16941, A2 => n17248, B1 => n13673, B2 => 
                           n16937, ZN => n1420);
   U16188 : OAI22_X1 port map( A1 => n16941, A2 => n17251, B1 => n13672, B2 => 
                           n16937, ZN => n1421);
   U16189 : OAI22_X1 port map( A1 => n16941, A2 => n17254, B1 => n13671, B2 => 
                           n16937, ZN => n1422);
   U16190 : OAI22_X1 port map( A1 => n16941, A2 => n17257, B1 => n13670, B2 => 
                           n16937, ZN => n1423);
   U16191 : OAI22_X1 port map( A1 => n16942, A2 => n17260, B1 => n13669, B2 => 
                           n16937, ZN => n1424);
   U16192 : OAI22_X1 port map( A1 => n16942, A2 => n17263, B1 => n13668, B2 => 
                           n16937, ZN => n1425);
   U16193 : OAI22_X1 port map( A1 => n16942, A2 => n17266, B1 => n13667, B2 => 
                           n16937, ZN => n1426);
   U16194 : OAI22_X1 port map( A1 => n16942, A2 => n17269, B1 => n13666, B2 => 
                           n16937, ZN => n1427);
   U16195 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_24_port, C1 => n16753,
                           C2 => n16414, A => n15924, ZN => n15912);
   U16196 : AOI21_X1 port map( B1 => n15925, B2 => n15926, A => n16750, ZN => 
                           n15924);
   U16197 : AOI221_X1 port map( B1 => n16735, B2 => n14892, C1 => n16732, C2 =>
                           n14908, A => n15928, ZN => n15925);
   U16198 : AOI221_X1 port map( B1 => n16745, B2 => n14884, C1 => n16742, C2 =>
                           n14900, A => n15927, ZN => n15926);
   U16199 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_25_port, C1 => n16753,
                           C2 => n16415, A => n15907, ZN => n15895);
   U16200 : AOI21_X1 port map( B1 => n15908, B2 => n15909, A => n16750, ZN => 
                           n15907);
   U16201 : AOI221_X1 port map( B1 => n16735, B2 => n14891, C1 => n16732, C2 =>
                           n14907, A => n15911, ZN => n15908);
   U16202 : AOI221_X1 port map( B1 => n16745, B2 => n14883, C1 => n16742, C2 =>
                           n14899, A => n15910, ZN => n15909);
   U16203 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_26_port, C1 => n16753,
                           C2 => n16416, A => n15890, ZN => n15878);
   U16204 : AOI21_X1 port map( B1 => n15891, B2 => n15892, A => n16750, ZN => 
                           n15890);
   U16205 : AOI221_X1 port map( B1 => n16735, B2 => n14890, C1 => n16732, C2 =>
                           n14906, A => n15894, ZN => n15891);
   U16206 : AOI221_X1 port map( B1 => n16745, B2 => n14882, C1 => n16742, C2 =>
                           n14898, A => n15893, ZN => n15892);
   U16207 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_27_port, C1 => n16753,
                           C2 => n16417, A => n15873, ZN => n15861);
   U16208 : AOI21_X1 port map( B1 => n15874, B2 => n15875, A => n16750, ZN => 
                           n15873);
   U16209 : AOI221_X1 port map( B1 => n16735, B2 => n14889, C1 => n16732, C2 =>
                           n14905, A => n15877, ZN => n15874);
   U16210 : AOI221_X1 port map( B1 => n16745, B2 => n14881, C1 => n16742, C2 =>
                           n14897, A => n15876, ZN => n15875);
   U16211 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_28_port, C1 => n16753,
                           C2 => n16418, A => n15856, ZN => n15844);
   U16212 : AOI21_X1 port map( B1 => n15857, B2 => n15858, A => n16750, ZN => 
                           n15856);
   U16213 : AOI221_X1 port map( B1 => n16735, B2 => n14888, C1 => n16732, C2 =>
                           n14904, A => n15860, ZN => n15857);
   U16214 : AOI221_X1 port map( B1 => n16745, B2 => n14880, C1 => n16742, C2 =>
                           n14896, A => n15859, ZN => n15858);
   U16215 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_29_port, C1 => n16753,
                           C2 => n16419, A => n15839, ZN => n15827);
   U16216 : AOI21_X1 port map( B1 => n15840, B2 => n15841, A => n16750, ZN => 
                           n15839);
   U16217 : AOI221_X1 port map( B1 => n16735, B2 => n14887, C1 => n16732, C2 =>
                           n14903, A => n15843, ZN => n15840);
   U16218 : AOI221_X1 port map( B1 => n16745, B2 => n14879, C1 => n16742, C2 =>
                           n14895, A => n15842, ZN => n15841);
   U16219 : AOI221_X1 port map( B1 => n16754, B2 => OUT2_30_port, C1 => n16753,
                           C2 => n16420, A => n15822, ZN => n15810);
   U16220 : AOI21_X1 port map( B1 => n15823, B2 => n15824, A => n16750, ZN => 
                           n15822);
   U16221 : AOI221_X1 port map( B1 => n16735, B2 => n14886, C1 => n16732, C2 =>
                           n14902, A => n15826, ZN => n15823);
   U16222 : AOI221_X1 port map( B1 => n16745, B2 => n14878, C1 => n16742, C2 =>
                           n14894, A => n15825, ZN => n15824);
   U16223 : AOI221_X1 port map( B1 => n16755, B2 => OUT2_31_port, C1 => n16753,
                           C2 => n16421, A => n15798, ZN => n15761);
   U16224 : AOI21_X1 port map( B1 => n15799, B2 => n15800, A => n16750, ZN => 
                           n15798);
   U16225 : AOI221_X1 port map( B1 => n16736, B2 => n14885, C1 => n16733, C2 =>
                           n14901, A => n15809, ZN => n15799);
   U16226 : AOI221_X1 port map( B1 => n16746, B2 => n14877, C1 => n16743, C2 =>
                           n14893, A => n15804, ZN => n15800);
   U16227 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_24_port, C1 => n16846,
                           C2 => n16414, A => n15343, ZN => n15331);
   U16228 : AOI21_X1 port map( B1 => n15344, B2 => n15345, A => n16843, ZN => 
                           n15343);
   U16229 : AOI221_X1 port map( B1 => n16828, B2 => n14892, C1 => n16825, C2 =>
                           n14908, A => n15347, ZN => n15344);
   U16230 : AOI221_X1 port map( B1 => n16838, B2 => n14884, C1 => n16835, C2 =>
                           n14900, A => n15346, ZN => n15345);
   U16231 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_25_port, C1 => n16846,
                           C2 => n16415, A => n15326, ZN => n15314);
   U16232 : AOI21_X1 port map( B1 => n15327, B2 => n15328, A => n16843, ZN => 
                           n15326);
   U16233 : AOI221_X1 port map( B1 => n16828, B2 => n14891, C1 => n16825, C2 =>
                           n14907, A => n15330, ZN => n15327);
   U16234 : AOI221_X1 port map( B1 => n16838, B2 => n14883, C1 => n16835, C2 =>
                           n14899, A => n15329, ZN => n15328);
   U16235 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_26_port, C1 => n16846,
                           C2 => n16416, A => n15309, ZN => n15297);
   U16236 : AOI21_X1 port map( B1 => n15310, B2 => n15311, A => n16843, ZN => 
                           n15309);
   U16237 : AOI221_X1 port map( B1 => n16828, B2 => n14890, C1 => n16825, C2 =>
                           n14906, A => n15313, ZN => n15310);
   U16238 : AOI221_X1 port map( B1 => n16838, B2 => n14882, C1 => n16835, C2 =>
                           n14898, A => n15312, ZN => n15311);
   U16239 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_27_port, C1 => n16846,
                           C2 => n16417, A => n15292, ZN => n15280);
   U16240 : AOI21_X1 port map( B1 => n15293, B2 => n15294, A => n16843, ZN => 
                           n15292);
   U16241 : AOI221_X1 port map( B1 => n16828, B2 => n14889, C1 => n16825, C2 =>
                           n14905, A => n15296, ZN => n15293);
   U16242 : AOI221_X1 port map( B1 => n16838, B2 => n14881, C1 => n16835, C2 =>
                           n14897, A => n15295, ZN => n15294);
   U16243 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_28_port, C1 => n16846,
                           C2 => n16418, A => n15275, ZN => n15263);
   U16244 : AOI21_X1 port map( B1 => n15276, B2 => n15277, A => n16843, ZN => 
                           n15275);
   U16245 : AOI221_X1 port map( B1 => n16828, B2 => n14888, C1 => n16825, C2 =>
                           n14904, A => n15279, ZN => n15276);
   U16246 : AOI221_X1 port map( B1 => n16838, B2 => n14880, C1 => n16835, C2 =>
                           n14896, A => n15278, ZN => n15277);
   U16247 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_29_port, C1 => n16846,
                           C2 => n16419, A => n15258, ZN => n15246);
   U16248 : AOI21_X1 port map( B1 => n15259, B2 => n15260, A => n16843, ZN => 
                           n15258);
   U16249 : AOI221_X1 port map( B1 => n16828, B2 => n14887, C1 => n16825, C2 =>
                           n14903, A => n15262, ZN => n15259);
   U16250 : AOI221_X1 port map( B1 => n16838, B2 => n14879, C1 => n16835, C2 =>
                           n14895, A => n15261, ZN => n15260);
   U16251 : AOI221_X1 port map( B1 => n16847, B2 => OUT1_30_port, C1 => n16846,
                           C2 => n16420, A => n15241, ZN => n15229);
   U16252 : AOI21_X1 port map( B1 => n15242, B2 => n15243, A => n16843, ZN => 
                           n15241);
   U16253 : AOI221_X1 port map( B1 => n16828, B2 => n14886, C1 => n16825, C2 =>
                           n14902, A => n15245, ZN => n15242);
   U16254 : AOI221_X1 port map( B1 => n16838, B2 => n14878, C1 => n16835, C2 =>
                           n14894, A => n15244, ZN => n15243);
   U16255 : AOI221_X1 port map( B1 => n16848, B2 => OUT1_31_port, C1 => n16846,
                           C2 => n16421, A => n15217, ZN => n15180);
   U16256 : AOI21_X1 port map( B1 => n15218, B2 => n15219, A => n16843, ZN => 
                           n15217);
   U16257 : AOI221_X1 port map( B1 => n16829, B2 => n14885, C1 => n16826, C2 =>
                           n14901, A => n15228, ZN => n15218);
   U16258 : AOI221_X1 port map( B1 => n16839, B2 => n14877, C1 => n16836, C2 =>
                           n14893, A => n15223, ZN => n15219);
   U16259 : NAND4_X1 port map( A1 => n16320, A2 => n16321, A3 => n16322, A4 => 
                           n16323, ZN => n1276);
   U16260 : AOI222_X1 port map( A1 => n16762, A2 => n16558, B1 => n16761, B2 =>
                           n16654, C1 => n16758, C2 => n16534, ZN => n16321);
   U16261 : NOR4_X1 port map( A1 => n16324, A2 => n16325, A3 => n16326, A4 => 
                           n16327, ZN => n16323);
   U16262 : AOI211_X1 port map( C1 => n16783, C2 => n16702, A => n16333, B => 
                           n16334, ZN => n16322);
   U16263 : NAND4_X1 port map( A1 => n16303, A2 => n16304, A3 => n16305, A4 => 
                           n16306, ZN => n1277);
   U16264 : AOI222_X1 port map( A1 => n16762, A2 => n16559, B1 => n16761, B2 =>
                           n16655, C1 => n16758, C2 => n16535, ZN => n16304);
   U16265 : NOR4_X1 port map( A1 => n16307, A2 => n16308, A3 => n16309, A4 => 
                           n16310, ZN => n16306);
   U16266 : AOI211_X1 port map( C1 => n16783, C2 => n16703, A => n16312, B => 
                           n16313, ZN => n16305);
   U16267 : NAND4_X1 port map( A1 => n16286, A2 => n16287, A3 => n16288, A4 => 
                           n16289, ZN => n1278);
   U16268 : AOI222_X1 port map( A1 => n16762, A2 => n16560, B1 => n16761, B2 =>
                           n16656, C1 => n16758, C2 => n16536, ZN => n16287);
   U16269 : NOR4_X1 port map( A1 => n16290, A2 => n16291, A3 => n16292, A4 => 
                           n16293, ZN => n16289);
   U16270 : AOI211_X1 port map( C1 => n16783, C2 => n16704, A => n16295, B => 
                           n16296, ZN => n16288);
   U16271 : NAND4_X1 port map( A1 => n16269, A2 => n16270, A3 => n16271, A4 => 
                           n16272, ZN => n1279);
   U16272 : AOI222_X1 port map( A1 => n16762, A2 => n16561, B1 => n16761, B2 =>
                           n16657, C1 => n16758, C2 => n16537, ZN => n16270);
   U16273 : NOR4_X1 port map( A1 => n16273, A2 => n16274, A3 => n16275, A4 => 
                           n16276, ZN => n16272);
   U16274 : AOI211_X1 port map( C1 => n16783, C2 => n16705, A => n16278, B => 
                           n16279, ZN => n16271);
   U16275 : NAND4_X1 port map( A1 => n16252, A2 => n16253, A3 => n16254, A4 => 
                           n16255, ZN => n1280);
   U16276 : AOI222_X1 port map( A1 => n16762, A2 => n16562, B1 => n16761, B2 =>
                           n16658, C1 => n16758, C2 => n16538, ZN => n16253);
   U16277 : NOR4_X1 port map( A1 => n16256, A2 => n16257, A3 => n16258, A4 => 
                           n16259, ZN => n16255);
   U16278 : AOI211_X1 port map( C1 => n16783, C2 => n16706, A => n16261, B => 
                           n16262, ZN => n16254);
   U16279 : NAND4_X1 port map( A1 => n16235, A2 => n16236, A3 => n16237, A4 => 
                           n16238, ZN => n1281);
   U16280 : AOI222_X1 port map( A1 => n16762, A2 => n16563, B1 => n16761, B2 =>
                           n16659, C1 => n16758, C2 => n16539, ZN => n16236);
   U16281 : NOR4_X1 port map( A1 => n16239, A2 => n16240, A3 => n16241, A4 => 
                           n16242, ZN => n16238);
   U16282 : AOI211_X1 port map( C1 => n16783, C2 => n16707, A => n16244, B => 
                           n16245, ZN => n16237);
   U16283 : NAND4_X1 port map( A1 => n16218, A2 => n16219, A3 => n16220, A4 => 
                           n16221, ZN => n1282);
   U16284 : AOI222_X1 port map( A1 => n16762, A2 => n16564, B1 => n16761, B2 =>
                           n16660, C1 => n16758, C2 => n16540, ZN => n16219);
   U16285 : NOR4_X1 port map( A1 => n16222, A2 => n16223, A3 => n16224, A4 => 
                           n16225, ZN => n16221);
   U16286 : AOI211_X1 port map( C1 => n16783, C2 => n16708, A => n16227, B => 
                           n16228, ZN => n16220);
   U16287 : NAND4_X1 port map( A1 => n16201, A2 => n16202, A3 => n16203, A4 => 
                           n16204, ZN => n1283);
   U16288 : AOI222_X1 port map( A1 => n16762, A2 => n16565, B1 => n16761, B2 =>
                           n16661, C1 => n16758, C2 => n16541, ZN => n16202);
   U16289 : NOR4_X1 port map( A1 => n16205, A2 => n16206, A3 => n16207, A4 => 
                           n16208, ZN => n16204);
   U16290 : AOI211_X1 port map( C1 => n16783, C2 => n16709, A => n16210, B => 
                           n16211, ZN => n16203);
   U16291 : NAND4_X1 port map( A1 => n16184, A2 => n16185, A3 => n16186, A4 => 
                           n16187, ZN => n1284);
   U16292 : AOI222_X1 port map( A1 => n16762, A2 => n16566, B1 => n16760, B2 =>
                           n16662, C1 => n16757, C2 => n16542, ZN => n16185);
   U16293 : NOR4_X1 port map( A1 => n16188, A2 => n16189, A3 => n16190, A4 => 
                           n16191, ZN => n16187);
   U16294 : AOI211_X1 port map( C1 => n16783, C2 => n16710, A => n16193, B => 
                           n16194, ZN => n16186);
   U16295 : NAND4_X1 port map( A1 => n16167, A2 => n16168, A3 => n16169, A4 => 
                           n16170, ZN => n1285);
   U16296 : AOI222_X1 port map( A1 => n16762, A2 => n16567, B1 => n16760, B2 =>
                           n16663, C1 => n16757, C2 => n16543, ZN => n16168);
   U16297 : NOR4_X1 port map( A1 => n16171, A2 => n16172, A3 => n16173, A4 => 
                           n16174, ZN => n16170);
   U16298 : AOI211_X1 port map( C1 => n16783, C2 => n16711, A => n16176, B => 
                           n16177, ZN => n16169);
   U16299 : NAND4_X1 port map( A1 => n16150, A2 => n16151, A3 => n16152, A4 => 
                           n16153, ZN => n1286);
   U16300 : AOI222_X1 port map( A1 => n16762, A2 => n16568, B1 => n16760, B2 =>
                           n16664, C1 => n16757, C2 => n16544, ZN => n16151);
   U16301 : NOR4_X1 port map( A1 => n16154, A2 => n16155, A3 => n16156, A4 => 
                           n16157, ZN => n16153);
   U16302 : AOI211_X1 port map( C1 => n16783, C2 => n16712, A => n16159, B => 
                           n16160, ZN => n16152);
   U16303 : NAND4_X1 port map( A1 => n16133, A2 => n16134, A3 => n16135, A4 => 
                           n16136, ZN => n1287);
   U16304 : AOI222_X1 port map( A1 => n16762, A2 => n16569, B1 => n16760, B2 =>
                           n16665, C1 => n16757, C2 => n16545, ZN => n16134);
   U16305 : NOR4_X1 port map( A1 => n16137, A2 => n16138, A3 => n16139, A4 => 
                           n16140, ZN => n16136);
   U16306 : AOI211_X1 port map( C1 => n16783, C2 => n16713, A => n16142, B => 
                           n16143, ZN => n16135);
   U16307 : NAND4_X1 port map( A1 => n16116, A2 => n16117, A3 => n16118, A4 => 
                           n16119, ZN => n1288);
   U16308 : AOI222_X1 port map( A1 => n16763, A2 => n16570, B1 => n16760, B2 =>
                           n16666, C1 => n16757, C2 => n16546, ZN => n16117);
   U16309 : NOR4_X1 port map( A1 => n16120, A2 => n16121, A3 => n16122, A4 => 
                           n16123, ZN => n16119);
   U16310 : AOI211_X1 port map( C1 => n16784, C2 => n16714, A => n16125, B => 
                           n16126, ZN => n16118);
   U16311 : NAND4_X1 port map( A1 => n16099, A2 => n16100, A3 => n16101, A4 => 
                           n16102, ZN => n1289);
   U16312 : AOI222_X1 port map( A1 => n16763, A2 => n16571, B1 => n16760, B2 =>
                           n16667, C1 => n16757, C2 => n16547, ZN => n16100);
   U16313 : NOR4_X1 port map( A1 => n16103, A2 => n16104, A3 => n16105, A4 => 
                           n16106, ZN => n16102);
   U16314 : AOI211_X1 port map( C1 => n16784, C2 => n16715, A => n16108, B => 
                           n16109, ZN => n16101);
   U16315 : NAND4_X1 port map( A1 => n16082, A2 => n16083, A3 => n16084, A4 => 
                           n16085, ZN => n1290);
   U16316 : AOI222_X1 port map( A1 => n16763, A2 => n16572, B1 => n16760, B2 =>
                           n16668, C1 => n16757, C2 => n16548, ZN => n16083);
   U16317 : NOR4_X1 port map( A1 => n16086, A2 => n16087, A3 => n16088, A4 => 
                           n16089, ZN => n16085);
   U16318 : AOI211_X1 port map( C1 => n16784, C2 => n16716, A => n16091, B => 
                           n16092, ZN => n16084);
   U16319 : NAND4_X1 port map( A1 => n16065, A2 => n16066, A3 => n16067, A4 => 
                           n16068, ZN => n1291);
   U16320 : AOI222_X1 port map( A1 => n16763, A2 => n16573, B1 => n16760, B2 =>
                           n16669, C1 => n16757, C2 => n16549, ZN => n16066);
   U16321 : NOR4_X1 port map( A1 => n16069, A2 => n16070, A3 => n16071, A4 => 
                           n16072, ZN => n16068);
   U16322 : AOI211_X1 port map( C1 => n16784, C2 => n16717, A => n16074, B => 
                           n16075, ZN => n16067);
   U16323 : NAND4_X1 port map( A1 => n16048, A2 => n16049, A3 => n16050, A4 => 
                           n16051, ZN => n1292);
   U16324 : AOI222_X1 port map( A1 => n16763, A2 => n16574, B1 => n16760, B2 =>
                           n16670, C1 => n16757, C2 => n16550, ZN => n16049);
   U16325 : NOR4_X1 port map( A1 => n16052, A2 => n16053, A3 => n16054, A4 => 
                           n16055, ZN => n16051);
   U16326 : AOI211_X1 port map( C1 => n16784, C2 => n16718, A => n16057, B => 
                           n16058, ZN => n16050);
   U16327 : NAND4_X1 port map( A1 => n16031, A2 => n16032, A3 => n16033, A4 => 
                           n16034, ZN => n1293);
   U16328 : AOI222_X1 port map( A1 => n16763, A2 => n16575, B1 => n16760, B2 =>
                           n16671, C1 => n16757, C2 => n16551, ZN => n16032);
   U16329 : NOR4_X1 port map( A1 => n16035, A2 => n16036, A3 => n16037, A4 => 
                           n16038, ZN => n16034);
   U16330 : AOI211_X1 port map( C1 => n16784, C2 => n16719, A => n16040, B => 
                           n16041, ZN => n16033);
   U16331 : NAND4_X1 port map( A1 => n16014, A2 => n16015, A3 => n16016, A4 => 
                           n16017, ZN => n1294);
   U16332 : AOI222_X1 port map( A1 => n16763, A2 => n16576, B1 => n16760, B2 =>
                           n16672, C1 => n16757, C2 => n16552, ZN => n16015);
   U16333 : NOR4_X1 port map( A1 => n16018, A2 => n16019, A3 => n16020, A4 => 
                           n16021, ZN => n16017);
   U16334 : AOI211_X1 port map( C1 => n16784, C2 => n16720, A => n16023, B => 
                           n16024, ZN => n16016);
   U16335 : NAND4_X1 port map( A1 => n15997, A2 => n15998, A3 => n15999, A4 => 
                           n16000, ZN => n1295);
   U16336 : AOI222_X1 port map( A1 => n16763, A2 => n16577, B1 => n16760, B2 =>
                           n16673, C1 => n16757, C2 => n16553, ZN => n15998);
   U16337 : NOR4_X1 port map( A1 => n16001, A2 => n16002, A3 => n16003, A4 => 
                           n16004, ZN => n16000);
   U16338 : AOI211_X1 port map( C1 => n16784, C2 => n16721, A => n16006, B => 
                           n16007, ZN => n15999);
   U16339 : NAND4_X1 port map( A1 => n15980, A2 => n15981, A3 => n15982, A4 => 
                           n15983, ZN => n1296);
   U16340 : AOI222_X1 port map( A1 => n16763, A2 => n16578, B1 => n16759, B2 =>
                           n16674, C1 => n16756, C2 => n16554, ZN => n15981);
   U16341 : NOR4_X1 port map( A1 => n15984, A2 => n15985, A3 => n15986, A4 => 
                           n15987, ZN => n15983);
   U16342 : AOI211_X1 port map( C1 => n16784, C2 => n16722, A => n15989, B => 
                           n15990, ZN => n15982);
   U16343 : NAND4_X1 port map( A1 => n15963, A2 => n15964, A3 => n15965, A4 => 
                           n15966, ZN => n1297);
   U16344 : AOI222_X1 port map( A1 => n16763, A2 => n16579, B1 => n16759, B2 =>
                           n16675, C1 => n16756, C2 => n16555, ZN => n15964);
   U16345 : NOR4_X1 port map( A1 => n15967, A2 => n15968, A3 => n15969, A4 => 
                           n15970, ZN => n15966);
   U16346 : AOI211_X1 port map( C1 => n16784, C2 => n16723, A => n15972, B => 
                           n15973, ZN => n15965);
   U16347 : NAND4_X1 port map( A1 => n15946, A2 => n15947, A3 => n15948, A4 => 
                           n15949, ZN => n1298);
   U16348 : AOI222_X1 port map( A1 => n16763, A2 => n16580, B1 => n16759, B2 =>
                           n16676, C1 => n16756, C2 => n16556, ZN => n15947);
   U16349 : NOR4_X1 port map( A1 => n15950, A2 => n15951, A3 => n15952, A4 => 
                           n15953, ZN => n15949);
   U16350 : AOI211_X1 port map( C1 => n16784, C2 => n16724, A => n15955, B => 
                           n15956, ZN => n15948);
   U16351 : NAND4_X1 port map( A1 => n15929, A2 => n15930, A3 => n15931, A4 => 
                           n15932, ZN => n1299);
   U16352 : AOI222_X1 port map( A1 => n16763, A2 => n16581, B1 => n16759, B2 =>
                           n16677, C1 => n16756, C2 => n16557, ZN => n15930);
   U16353 : NOR4_X1 port map( A1 => n15933, A2 => n15934, A3 => n15935, A4 => 
                           n15936, ZN => n15932);
   U16354 : AOI211_X1 port map( C1 => n16784, C2 => n16725, A => n15938, B => 
                           n15939, ZN => n15931);
   U16355 : NAND4_X1 port map( A1 => n15912, A2 => n15913, A3 => n15914, A4 => 
                           n15915, ZN => n1300);
   U16356 : AOI222_X1 port map( A1 => n16764, A2 => n16430, B1 => n16759, B2 =>
                           n16366, C1 => n16756, C2 => n16422, ZN => n15913);
   U16357 : NOR4_X1 port map( A1 => n15916, A2 => n15917, A3 => n15918, A4 => 
                           n15919, ZN => n15915);
   U16358 : AOI211_X1 port map( C1 => n16785, C2 => n16382, A => n15921, B => 
                           n15922, ZN => n15914);
   U16359 : NAND4_X1 port map( A1 => n15895, A2 => n15896, A3 => n15897, A4 => 
                           n15898, ZN => n1301);
   U16360 : AOI222_X1 port map( A1 => n16764, A2 => n16431, B1 => n16759, B2 =>
                           n16367, C1 => n16756, C2 => n16423, ZN => n15896);
   U16361 : NOR4_X1 port map( A1 => n15899, A2 => n15900, A3 => n15901, A4 => 
                           n15902, ZN => n15898);
   U16362 : AOI211_X1 port map( C1 => n16785, C2 => n16383, A => n15904, B => 
                           n15905, ZN => n15897);
   U16363 : NAND4_X1 port map( A1 => n15878, A2 => n15879, A3 => n15880, A4 => 
                           n15881, ZN => n1302);
   U16364 : AOI222_X1 port map( A1 => n16764, A2 => n16432, B1 => n16759, B2 =>
                           n16368, C1 => n16756, C2 => n16424, ZN => n15879);
   U16365 : NOR4_X1 port map( A1 => n15882, A2 => n15883, A3 => n15884, A4 => 
                           n15885, ZN => n15881);
   U16366 : AOI211_X1 port map( C1 => n16785, C2 => n16384, A => n15887, B => 
                           n15888, ZN => n15880);
   U16367 : NAND4_X1 port map( A1 => n15861, A2 => n15862, A3 => n15863, A4 => 
                           n15864, ZN => n1303);
   U16368 : AOI222_X1 port map( A1 => n16764, A2 => n16433, B1 => n16759, B2 =>
                           n16369, C1 => n16756, C2 => n16425, ZN => n15862);
   U16369 : NOR4_X1 port map( A1 => n15865, A2 => n15866, A3 => n15867, A4 => 
                           n15868, ZN => n15864);
   U16370 : AOI211_X1 port map( C1 => n16785, C2 => n16385, A => n15870, B => 
                           n15871, ZN => n15863);
   U16371 : NAND4_X1 port map( A1 => n15844, A2 => n15845, A3 => n15846, A4 => 
                           n15847, ZN => n1304);
   U16372 : AOI222_X1 port map( A1 => n16764, A2 => n16434, B1 => n16759, B2 =>
                           n16370, C1 => n16756, C2 => n16426, ZN => n15845);
   U16373 : NOR4_X1 port map( A1 => n15848, A2 => n15849, A3 => n15850, A4 => 
                           n15851, ZN => n15847);
   U16374 : AOI211_X1 port map( C1 => n16785, C2 => n16386, A => n15853, B => 
                           n15854, ZN => n15846);
   U16375 : NAND4_X1 port map( A1 => n15827, A2 => n15828, A3 => n15829, A4 => 
                           n15830, ZN => n1305);
   U16376 : AOI222_X1 port map( A1 => n16764, A2 => n16435, B1 => n16759, B2 =>
                           n16371, C1 => n16756, C2 => n16427, ZN => n15828);
   U16377 : NOR4_X1 port map( A1 => n15831, A2 => n15832, A3 => n15833, A4 => 
                           n15834, ZN => n15830);
   U16378 : AOI211_X1 port map( C1 => n16785, C2 => n16387, A => n15836, B => 
                           n15837, ZN => n15829);
   U16379 : NAND4_X1 port map( A1 => n15810, A2 => n15811, A3 => n15812, A4 => 
                           n15813, ZN => n1306);
   U16380 : AOI222_X1 port map( A1 => n16764, A2 => n16436, B1 => n16759, B2 =>
                           n16372, C1 => n16756, C2 => n16428, ZN => n15811);
   U16381 : NOR4_X1 port map( A1 => n15814, A2 => n15815, A3 => n15816, A4 => 
                           n15817, ZN => n15813);
   U16382 : AOI211_X1 port map( C1 => n16785, C2 => n16388, A => n15819, B => 
                           n15820, ZN => n15812);
   U16383 : NAND4_X1 port map( A1 => n15761, A2 => n15762, A3 => n15763, A4 => 
                           n15764, ZN => n1307);
   U16384 : AOI222_X1 port map( A1 => n16764, A2 => n16437, B1 => n16759, B2 =>
                           n16373, C1 => n16756, C2 => n16429, ZN => n15762);
   U16385 : NOR4_X1 port map( A1 => n15765, A2 => n15766, A3 => n15767, A4 => 
                           n15768, ZN => n15764);
   U16386 : AOI211_X1 port map( C1 => n16785, C2 => n16389, A => n15784, B => 
                           n15785, ZN => n15763);
   U16387 : NAND4_X1 port map( A1 => n15739, A2 => n15740, A3 => n15741, A4 => 
                           n15742, ZN => n1308);
   U16388 : AOI222_X1 port map( A1 => n16855, A2 => n16558, B1 => n16854, B2 =>
                           n16654, C1 => n16851, C2 => n16534, ZN => n15740);
   U16389 : NOR4_X1 port map( A1 => n15743, A2 => n15744, A3 => n15745, A4 => 
                           n15746, ZN => n15742);
   U16390 : AOI211_X1 port map( C1 => n16876, C2 => n16702, A => n15752, B => 
                           n15753, ZN => n15741);
   U16391 : NAND4_X1 port map( A1 => n15722, A2 => n15723, A3 => n15724, A4 => 
                           n15725, ZN => n1309);
   U16392 : AOI222_X1 port map( A1 => n16855, A2 => n16559, B1 => n16854, B2 =>
                           n16655, C1 => n16851, C2 => n16535, ZN => n15723);
   U16393 : NOR4_X1 port map( A1 => n15726, A2 => n15727, A3 => n15728, A4 => 
                           n15729, ZN => n15725);
   U16394 : AOI211_X1 port map( C1 => n16876, C2 => n16703, A => n15731, B => 
                           n15732, ZN => n15724);
   U16395 : NAND4_X1 port map( A1 => n15705, A2 => n15706, A3 => n15707, A4 => 
                           n15708, ZN => n1310);
   U16396 : AOI222_X1 port map( A1 => n16855, A2 => n16560, B1 => n16854, B2 =>
                           n16656, C1 => n16851, C2 => n16536, ZN => n15706);
   U16397 : NOR4_X1 port map( A1 => n15709, A2 => n15710, A3 => n15711, A4 => 
                           n15712, ZN => n15708);
   U16398 : AOI211_X1 port map( C1 => n16876, C2 => n16704, A => n15714, B => 
                           n15715, ZN => n15707);
   U16399 : NAND4_X1 port map( A1 => n15688, A2 => n15689, A3 => n15690, A4 => 
                           n15691, ZN => n1311);
   U16400 : AOI222_X1 port map( A1 => n16855, A2 => n16561, B1 => n16854, B2 =>
                           n16657, C1 => n16851, C2 => n16537, ZN => n15689);
   U16401 : NOR4_X1 port map( A1 => n15692, A2 => n15693, A3 => n15694, A4 => 
                           n15695, ZN => n15691);
   U16402 : AOI211_X1 port map( C1 => n16876, C2 => n16705, A => n15697, B => 
                           n15698, ZN => n15690);
   U16403 : NAND4_X1 port map( A1 => n15671, A2 => n15672, A3 => n15673, A4 => 
                           n15674, ZN => n1312);
   U16404 : AOI222_X1 port map( A1 => n16855, A2 => n16562, B1 => n16854, B2 =>
                           n16658, C1 => n16851, C2 => n16538, ZN => n15672);
   U16405 : NOR4_X1 port map( A1 => n15675, A2 => n15676, A3 => n15677, A4 => 
                           n15678, ZN => n15674);
   U16406 : AOI211_X1 port map( C1 => n16876, C2 => n16706, A => n15680, B => 
                           n15681, ZN => n15673);
   U16407 : NAND4_X1 port map( A1 => n15654, A2 => n15655, A3 => n15656, A4 => 
                           n15657, ZN => n1313);
   U16408 : AOI222_X1 port map( A1 => n16855, A2 => n16563, B1 => n16854, B2 =>
                           n16659, C1 => n16851, C2 => n16539, ZN => n15655);
   U16409 : NOR4_X1 port map( A1 => n15658, A2 => n15659, A3 => n15660, A4 => 
                           n15661, ZN => n15657);
   U16410 : AOI211_X1 port map( C1 => n16876, C2 => n16707, A => n15663, B => 
                           n15664, ZN => n15656);
   U16411 : NAND4_X1 port map( A1 => n15637, A2 => n15638, A3 => n15639, A4 => 
                           n15640, ZN => n1314);
   U16412 : AOI222_X1 port map( A1 => n16855, A2 => n16564, B1 => n16854, B2 =>
                           n16660, C1 => n16851, C2 => n16540, ZN => n15638);
   U16413 : NOR4_X1 port map( A1 => n15641, A2 => n15642, A3 => n15643, A4 => 
                           n15644, ZN => n15640);
   U16414 : AOI211_X1 port map( C1 => n16876, C2 => n16708, A => n15646, B => 
                           n15647, ZN => n15639);
   U16415 : NAND4_X1 port map( A1 => n15620, A2 => n15621, A3 => n15622, A4 => 
                           n15623, ZN => n1315);
   U16416 : AOI222_X1 port map( A1 => n16855, A2 => n16565, B1 => n16854, B2 =>
                           n16661, C1 => n16851, C2 => n16541, ZN => n15621);
   U16417 : NOR4_X1 port map( A1 => n15624, A2 => n15625, A3 => n15626, A4 => 
                           n15627, ZN => n15623);
   U16418 : AOI211_X1 port map( C1 => n16876, C2 => n16709, A => n15629, B => 
                           n15630, ZN => n15622);
   U16419 : NAND4_X1 port map( A1 => n15603, A2 => n15604, A3 => n15605, A4 => 
                           n15606, ZN => n1316);
   U16420 : AOI222_X1 port map( A1 => n16855, A2 => n16566, B1 => n16853, B2 =>
                           n16662, C1 => n16850, C2 => n16542, ZN => n15604);
   U16421 : NOR4_X1 port map( A1 => n15607, A2 => n15608, A3 => n15609, A4 => 
                           n15610, ZN => n15606);
   U16422 : AOI211_X1 port map( C1 => n16876, C2 => n16710, A => n15612, B => 
                           n15613, ZN => n15605);
   U16423 : NAND4_X1 port map( A1 => n15586, A2 => n15587, A3 => n15588, A4 => 
                           n15589, ZN => n1317);
   U16424 : AOI222_X1 port map( A1 => n16855, A2 => n16567, B1 => n16853, B2 =>
                           n16663, C1 => n16850, C2 => n16543, ZN => n15587);
   U16425 : NOR4_X1 port map( A1 => n15590, A2 => n15591, A3 => n15592, A4 => 
                           n15593, ZN => n15589);
   U16426 : AOI211_X1 port map( C1 => n16876, C2 => n16711, A => n15595, B => 
                           n15596, ZN => n15588);
   U16427 : NAND4_X1 port map( A1 => n15569, A2 => n15570, A3 => n15571, A4 => 
                           n15572, ZN => n1318);
   U16428 : AOI222_X1 port map( A1 => n16855, A2 => n16568, B1 => n16853, B2 =>
                           n16664, C1 => n16850, C2 => n16544, ZN => n15570);
   U16429 : NOR4_X1 port map( A1 => n15573, A2 => n15574, A3 => n15575, A4 => 
                           n15576, ZN => n15572);
   U16430 : AOI211_X1 port map( C1 => n16876, C2 => n16712, A => n15578, B => 
                           n15579, ZN => n15571);
   U16431 : NAND4_X1 port map( A1 => n15552, A2 => n15553, A3 => n15554, A4 => 
                           n15555, ZN => n1319);
   U16432 : AOI222_X1 port map( A1 => n16855, A2 => n16569, B1 => n16853, B2 =>
                           n16665, C1 => n16850, C2 => n16545, ZN => n15553);
   U16433 : NOR4_X1 port map( A1 => n15556, A2 => n15557, A3 => n15558, A4 => 
                           n15559, ZN => n15555);
   U16434 : AOI211_X1 port map( C1 => n16876, C2 => n16713, A => n15561, B => 
                           n15562, ZN => n15554);
   U16435 : NAND4_X1 port map( A1 => n15535, A2 => n15536, A3 => n15537, A4 => 
                           n15538, ZN => n1320);
   U16436 : AOI222_X1 port map( A1 => n16856, A2 => n16570, B1 => n16853, B2 =>
                           n16666, C1 => n16850, C2 => n16546, ZN => n15536);
   U16437 : NOR4_X1 port map( A1 => n15539, A2 => n15540, A3 => n15541, A4 => 
                           n15542, ZN => n15538);
   U16438 : AOI211_X1 port map( C1 => n16877, C2 => n16714, A => n15544, B => 
                           n15545, ZN => n15537);
   U16439 : NAND4_X1 port map( A1 => n15518, A2 => n15519, A3 => n15520, A4 => 
                           n15521, ZN => n1321);
   U16440 : AOI222_X1 port map( A1 => n16856, A2 => n16571, B1 => n16853, B2 =>
                           n16667, C1 => n16850, C2 => n16547, ZN => n15519);
   U16441 : NOR4_X1 port map( A1 => n15522, A2 => n15523, A3 => n15524, A4 => 
                           n15525, ZN => n15521);
   U16442 : AOI211_X1 port map( C1 => n16877, C2 => n16715, A => n15527, B => 
                           n15528, ZN => n15520);
   U16443 : NAND4_X1 port map( A1 => n15501, A2 => n15502, A3 => n15503, A4 => 
                           n15504, ZN => n1322);
   U16444 : AOI222_X1 port map( A1 => n16856, A2 => n16572, B1 => n16853, B2 =>
                           n16668, C1 => n16850, C2 => n16548, ZN => n15502);
   U16445 : NOR4_X1 port map( A1 => n15505, A2 => n15506, A3 => n15507, A4 => 
                           n15508, ZN => n15504);
   U16446 : AOI211_X1 port map( C1 => n16877, C2 => n16716, A => n15510, B => 
                           n15511, ZN => n15503);
   U16447 : NAND4_X1 port map( A1 => n15484, A2 => n15485, A3 => n15486, A4 => 
                           n15487, ZN => n1323);
   U16448 : AOI222_X1 port map( A1 => n16856, A2 => n16573, B1 => n16853, B2 =>
                           n16669, C1 => n16850, C2 => n16549, ZN => n15485);
   U16449 : NOR4_X1 port map( A1 => n15488, A2 => n15489, A3 => n15490, A4 => 
                           n15491, ZN => n15487);
   U16450 : AOI211_X1 port map( C1 => n16877, C2 => n16717, A => n15493, B => 
                           n15494, ZN => n15486);
   U16451 : NAND4_X1 port map( A1 => n15467, A2 => n15468, A3 => n15469, A4 => 
                           n15470, ZN => n1324);
   U16452 : AOI222_X1 port map( A1 => n16856, A2 => n16574, B1 => n16853, B2 =>
                           n16670, C1 => n16850, C2 => n16550, ZN => n15468);
   U16453 : NOR4_X1 port map( A1 => n15471, A2 => n15472, A3 => n15473, A4 => 
                           n15474, ZN => n15470);
   U16454 : AOI211_X1 port map( C1 => n16877, C2 => n16718, A => n15476, B => 
                           n15477, ZN => n15469);
   U16455 : NAND4_X1 port map( A1 => n15450, A2 => n15451, A3 => n15452, A4 => 
                           n15453, ZN => n1325);
   U16456 : AOI222_X1 port map( A1 => n16856, A2 => n16575, B1 => n16853, B2 =>
                           n16671, C1 => n16850, C2 => n16551, ZN => n15451);
   U16457 : NOR4_X1 port map( A1 => n15454, A2 => n15455, A3 => n15456, A4 => 
                           n15457, ZN => n15453);
   U16458 : AOI211_X1 port map( C1 => n16877, C2 => n16719, A => n15459, B => 
                           n15460, ZN => n15452);
   U16459 : NAND4_X1 port map( A1 => n15433, A2 => n15434, A3 => n15435, A4 => 
                           n15436, ZN => n1326);
   U16460 : AOI222_X1 port map( A1 => n16856, A2 => n16576, B1 => n16853, B2 =>
                           n16672, C1 => n16850, C2 => n16552, ZN => n15434);
   U16461 : NOR4_X1 port map( A1 => n15437, A2 => n15438, A3 => n15439, A4 => 
                           n15440, ZN => n15436);
   U16462 : AOI211_X1 port map( C1 => n16877, C2 => n16720, A => n15442, B => 
                           n15443, ZN => n15435);
   U16463 : NAND4_X1 port map( A1 => n15416, A2 => n15417, A3 => n15418, A4 => 
                           n15419, ZN => n1327);
   U16464 : AOI222_X1 port map( A1 => n16856, A2 => n16577, B1 => n16853, B2 =>
                           n16673, C1 => n16850, C2 => n16553, ZN => n15417);
   U16465 : NOR4_X1 port map( A1 => n15420, A2 => n15421, A3 => n15422, A4 => 
                           n15423, ZN => n15419);
   U16466 : AOI211_X1 port map( C1 => n16877, C2 => n16721, A => n15425, B => 
                           n15426, ZN => n15418);
   U16467 : NAND4_X1 port map( A1 => n15399, A2 => n15400, A3 => n15401, A4 => 
                           n15402, ZN => n1328);
   U16468 : AOI222_X1 port map( A1 => n16856, A2 => n16578, B1 => n16852, B2 =>
                           n16674, C1 => n16849, C2 => n16554, ZN => n15400);
   U16469 : NOR4_X1 port map( A1 => n15403, A2 => n15404, A3 => n15405, A4 => 
                           n15406, ZN => n15402);
   U16470 : AOI211_X1 port map( C1 => n16877, C2 => n16722, A => n15408, B => 
                           n15409, ZN => n15401);
   U16471 : NAND4_X1 port map( A1 => n15382, A2 => n15383, A3 => n15384, A4 => 
                           n15385, ZN => n1329);
   U16472 : AOI222_X1 port map( A1 => n16856, A2 => n16579, B1 => n16852, B2 =>
                           n16675, C1 => n16849, C2 => n16555, ZN => n15383);
   U16473 : NOR4_X1 port map( A1 => n15386, A2 => n15387, A3 => n15388, A4 => 
                           n15389, ZN => n15385);
   U16474 : AOI211_X1 port map( C1 => n16877, C2 => n16723, A => n15391, B => 
                           n15392, ZN => n15384);
   U16475 : NAND4_X1 port map( A1 => n15365, A2 => n15366, A3 => n15367, A4 => 
                           n15368, ZN => n1330);
   U16476 : AOI222_X1 port map( A1 => n16856, A2 => n16580, B1 => n16852, B2 =>
                           n16676, C1 => n16849, C2 => n16556, ZN => n15366);
   U16477 : NOR4_X1 port map( A1 => n15369, A2 => n15370, A3 => n15371, A4 => 
                           n15372, ZN => n15368);
   U16478 : AOI211_X1 port map( C1 => n16877, C2 => n16724, A => n15374, B => 
                           n15375, ZN => n15367);
   U16479 : NAND4_X1 port map( A1 => n15348, A2 => n15349, A3 => n15350, A4 => 
                           n15351, ZN => n1331);
   U16480 : AOI222_X1 port map( A1 => n16856, A2 => n16581, B1 => n16852, B2 =>
                           n16677, C1 => n16849, C2 => n16557, ZN => n15349);
   U16481 : NOR4_X1 port map( A1 => n15352, A2 => n15353, A3 => n15354, A4 => 
                           n15355, ZN => n15351);
   U16482 : AOI211_X1 port map( C1 => n16877, C2 => n16725, A => n15357, B => 
                           n15358, ZN => n15350);
   U16483 : NAND4_X1 port map( A1 => n15331, A2 => n15332, A3 => n15333, A4 => 
                           n15334, ZN => n1332);
   U16484 : AOI222_X1 port map( A1 => n16857, A2 => n16430, B1 => n16852, B2 =>
                           n16366, C1 => n16849, C2 => n16422, ZN => n15332);
   U16485 : NOR4_X1 port map( A1 => n15335, A2 => n15336, A3 => n15337, A4 => 
                           n15338, ZN => n15334);
   U16486 : AOI211_X1 port map( C1 => n16878, C2 => n16382, A => n15340, B => 
                           n15341, ZN => n15333);
   U16487 : NAND4_X1 port map( A1 => n15314, A2 => n15315, A3 => n15316, A4 => 
                           n15317, ZN => n1333);
   U16488 : AOI222_X1 port map( A1 => n16857, A2 => n16431, B1 => n16852, B2 =>
                           n16367, C1 => n16849, C2 => n16423, ZN => n15315);
   U16489 : NOR4_X1 port map( A1 => n15318, A2 => n15319, A3 => n15320, A4 => 
                           n15321, ZN => n15317);
   U16490 : AOI211_X1 port map( C1 => n16878, C2 => n16383, A => n15323, B => 
                           n15324, ZN => n15316);
   U16491 : NAND4_X1 port map( A1 => n15297, A2 => n15298, A3 => n15299, A4 => 
                           n15300, ZN => n1334);
   U16492 : AOI222_X1 port map( A1 => n16857, A2 => n16432, B1 => n16852, B2 =>
                           n16368, C1 => n16849, C2 => n16424, ZN => n15298);
   U16493 : NOR4_X1 port map( A1 => n15301, A2 => n15302, A3 => n15303, A4 => 
                           n15304, ZN => n15300);
   U16494 : AOI211_X1 port map( C1 => n16878, C2 => n16384, A => n15306, B => 
                           n15307, ZN => n15299);
   U16495 : NAND4_X1 port map( A1 => n15280, A2 => n15281, A3 => n15282, A4 => 
                           n15283, ZN => n1335);
   U16496 : AOI222_X1 port map( A1 => n16857, A2 => n16433, B1 => n16852, B2 =>
                           n16369, C1 => n16849, C2 => n16425, ZN => n15281);
   U16497 : NOR4_X1 port map( A1 => n15284, A2 => n15285, A3 => n15286, A4 => 
                           n15287, ZN => n15283);
   U16498 : AOI211_X1 port map( C1 => n16878, C2 => n16385, A => n15289, B => 
                           n15290, ZN => n15282);
   U16499 : NAND4_X1 port map( A1 => n15263, A2 => n15264, A3 => n15265, A4 => 
                           n15266, ZN => n1336);
   U16500 : AOI222_X1 port map( A1 => n16857, A2 => n16434, B1 => n16852, B2 =>
                           n16370, C1 => n16849, C2 => n16426, ZN => n15264);
   U16501 : NOR4_X1 port map( A1 => n15267, A2 => n15268, A3 => n15269, A4 => 
                           n15270, ZN => n15266);
   U16502 : AOI211_X1 port map( C1 => n16878, C2 => n16386, A => n15272, B => 
                           n15273, ZN => n15265);
   U16503 : NAND4_X1 port map( A1 => n15246, A2 => n15247, A3 => n15248, A4 => 
                           n15249, ZN => n1337);
   U16504 : AOI222_X1 port map( A1 => n16857, A2 => n16435, B1 => n16852, B2 =>
                           n16371, C1 => n16849, C2 => n16427, ZN => n15247);
   U16505 : NOR4_X1 port map( A1 => n15250, A2 => n15251, A3 => n15252, A4 => 
                           n15253, ZN => n15249);
   U16506 : AOI211_X1 port map( C1 => n16878, C2 => n16387, A => n15255, B => 
                           n15256, ZN => n15248);
   U16507 : NAND4_X1 port map( A1 => n15229, A2 => n15230, A3 => n15231, A4 => 
                           n15232, ZN => n1338);
   U16508 : AOI222_X1 port map( A1 => n16857, A2 => n16436, B1 => n16852, B2 =>
                           n16372, C1 => n16849, C2 => n16428, ZN => n15230);
   U16509 : NOR4_X1 port map( A1 => n15233, A2 => n15234, A3 => n15235, A4 => 
                           n15236, ZN => n15232);
   U16510 : AOI211_X1 port map( C1 => n16878, C2 => n16388, A => n15238, B => 
                           n15239, ZN => n15231);
   U16511 : NAND4_X1 port map( A1 => n15180, A2 => n15181, A3 => n15182, A4 => 
                           n15183, ZN => n1339);
   U16512 : AOI222_X1 port map( A1 => n16857, A2 => n16437, B1 => n16852, B2 =>
                           n16373, C1 => n16849, C2 => n16429, ZN => n15181);
   U16513 : NOR4_X1 port map( A1 => n15184, A2 => n15185, A3 => n15186, A4 => 
                           n15187, ZN => n15183);
   U16514 : AOI211_X1 port map( C1 => n16878, C2 => n16389, A => n15203, B => 
                           n15204, ZN => n15182);
   U16515 : OAI22_X1 port map( A1 => n17109, A2 => n17198, B1 => n17108, B2 => 
                           n14749, ZN => n2012);
   U16516 : OAI22_X1 port map( A1 => n17109, A2 => n17201, B1 => n17108, B2 => 
                           n14748, ZN => n2013);
   U16517 : OAI22_X1 port map( A1 => n17109, A2 => n17204, B1 => n17108, B2 => 
                           n14747, ZN => n2014);
   U16518 : OAI22_X1 port map( A1 => n17109, A2 => n17207, B1 => n17108, B2 => 
                           n14746, ZN => n2015);
   U16519 : OAI22_X1 port map( A1 => n17109, A2 => n17210, B1 => n17108, B2 => 
                           n14745, ZN => n2016);
   U16520 : OAI22_X1 port map( A1 => n17110, A2 => n17213, B1 => n17108, B2 => 
                           n14744, ZN => n2017);
   U16521 : OAI22_X1 port map( A1 => n17110, A2 => n17216, B1 => n17108, B2 => 
                           n14743, ZN => n2018);
   U16522 : OAI22_X1 port map( A1 => n17110, A2 => n17219, B1 => n17108, B2 => 
                           n14742, ZN => n2019);
   U16523 : OAI22_X1 port map( A1 => n17110, A2 => n17222, B1 => n17108, B2 => 
                           n14741, ZN => n2020);
   U16524 : OAI22_X1 port map( A1 => n17110, A2 => n17225, B1 => n17108, B2 => 
                           n14740, ZN => n2021);
   U16525 : OAI22_X1 port map( A1 => n17111, A2 => n17228, B1 => n17108, B2 => 
                           n14739, ZN => n2022);
   U16526 : OAI22_X1 port map( A1 => n17111, A2 => n17231, B1 => n17108, B2 => 
                           n14738, ZN => n2023);
   U16527 : OAI22_X1 port map( A1 => n17111, A2 => n17234, B1 => n15152, B2 => 
                           n14737, ZN => n2024);
   U16528 : OAI22_X1 port map( A1 => n17111, A2 => n17237, B1 => n15152, B2 => 
                           n14736, ZN => n2025);
   U16529 : OAI22_X1 port map( A1 => n17111, A2 => n17240, B1 => n15152, B2 => 
                           n14735, ZN => n2026);
   U16530 : OAI22_X1 port map( A1 => n17112, A2 => n17243, B1 => n17108, B2 => 
                           n14734, ZN => n2027);
   U16531 : OAI22_X1 port map( A1 => n17112, A2 => n17246, B1 => n17108, B2 => 
                           n14733, ZN => n2028);
   U16532 : OAI22_X1 port map( A1 => n17112, A2 => n17249, B1 => n17108, B2 => 
                           n14732, ZN => n2029);
   U16533 : OAI22_X1 port map( A1 => n17112, A2 => n17252, B1 => n17108, B2 => 
                           n14731, ZN => n2030);
   U16534 : OAI22_X1 port map( A1 => n17112, A2 => n17255, B1 => n17108, B2 => 
                           n14730, ZN => n2031);
   U16535 : OAI22_X1 port map( A1 => n17113, A2 => n17258, B1 => n17108, B2 => 
                           n14729, ZN => n2032);
   U16536 : OAI22_X1 port map( A1 => n17113, A2 => n17261, B1 => n17108, B2 => 
                           n14728, ZN => n2033);
   U16537 : OAI22_X1 port map( A1 => n17113, A2 => n17264, B1 => n17108, B2 => 
                           n14727, ZN => n2034);
   U16538 : OAI22_X1 port map( A1 => n17113, A2 => n17267, B1 => n17108, B2 => 
                           n14726, ZN => n2035);
   U16539 : NOR3_X1 port map( A1 => n14460, A2 => ADD_RD2(2), A3 => n14459, ZN 
                           => n16328);
   U16540 : NOR3_X1 port map( A1 => n14453, A2 => ADD_RD1(2), A3 => n14452, ZN 
                           => n15747);
   U16541 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(3), A3 => n14459,
                           ZN => n16335);
   U16542 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(3), A3 => n14452,
                           ZN => n15754);
   U16543 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n15142);
   U16544 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n14447, ZN => n15140);
   U16545 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n14446, ZN => n15138);
   U16546 : AND3_X1 port map( A1 => n16726, A2 => n14461, A3 => ADD_RD2(0), ZN 
                           => n16329);
   U16547 : AND3_X1 port map( A1 => n16727, A2 => n14454, A3 => ADD_RD1(0), ZN 
                           => n15748);
   U16548 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(4), A3 => n14460,
                           ZN => n15807);
   U16549 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(4), A3 => n14453,
                           ZN => n15226);
   U16550 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(2), ZN => n15808);
   U16551 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(2), ZN => n15227);
   U16552 : INV_X1 port map( A => RESET, ZN => n14442);
   U16553 : AND3_X1 port map( A1 => ENABLE, A2 => n17320, A3 => RD2, ZN => 
                           n16726);
   U16554 : AND3_X1 port map( A1 => ENABLE, A2 => n17320, A3 => RD1, ZN => 
                           n16727);
   U16555 : AND3_X1 port map( A1 => n14460, A2 => n14459, A3 => ADD_RD2(2), ZN 
                           => n15803);
   U16556 : AND3_X1 port map( A1 => n14453, A2 => n14452, A3 => ADD_RD1(2), ZN 
                           => n15222);
   U16557 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n14459, A3 => ADD_RD2(3),
                           ZN => n15802);
   U16558 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n14452, A3 => ADD_RD1(3),
                           ZN => n15221);
   U16559 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n17316, ZN => n15127);
   U16560 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n17316, ZN => n15125);
   U16561 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n17316, ZN => n15124);
   U16562 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n17316, ZN => n15123);
   U16563 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n17316, ZN => n15122);
   U16564 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n17316, ZN => n15121);
   U16565 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n17316, ZN => n15120);
   U16566 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n17316, ZN => n15119);
   U16567 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n17316, ZN => n15118);
   U16568 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n17316, ZN => n15117);
   U16569 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n17316, ZN => n15116);
   U16570 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n17316, ZN => n15115);
   U16571 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n17315, ZN => n15114);
   U16572 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n17315, ZN => n15113);
   U16573 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n17315, ZN => n15112);
   U16574 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n17315, ZN => n15111);
   U16575 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n17315, ZN => n15110);
   U16576 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n17315, ZN => n15109);
   U16577 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n17315, ZN => n15108);
   U16578 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n17315, ZN => n15107);
   U16579 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n17315, ZN => n15106);
   U16580 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n17315, ZN => n15105);
   U16581 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n17315, ZN => n15104);
   U16582 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n17315, ZN => n15102);
   U16583 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n17317, ZN => n15134);
   U16584 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n17317, ZN => n15133);
   U16585 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n17317, ZN => n15132);
   U16586 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n17317, ZN => n15131);
   U16587 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n17317, ZN => n15130);
   U16588 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n17317, ZN => n15129);
   U16589 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n17317, ZN => n15128);
   U16590 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n17317, ZN => n15126);
   U16591 : INV_X1 port map( A => ADD_RD2(4), ZN => n14459);
   U16592 : INV_X1 port map( A => ADD_RD1(4), ZN => n14452);
   U16593 : INV_X1 port map( A => ADD_RD2(3), ZN => n14460);
   U16594 : INV_X1 port map( A => ADD_RD1(3), ZN => n14453);
   U16595 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n14460, A3 => ADD_RD2(4),
                           ZN => n16728);
   U16596 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n14453, A3 => ADD_RD1(4),
                           ZN => n16729);
   U16597 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n15164);
   U16598 : AND3_X1 port map( A1 => ENABLE, A2 => n14443, A3 => WR, ZN => 
                           n15143);
   U16599 : INV_X1 port map( A => ADD_WR(4), ZN => n14443);
   U16600 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(4), ZN => n16730);
   U16601 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(4), ZN => n16731);
   U16602 : INV_X1 port map( A => ADD_WR(3), ZN => n14444);
   U16603 : INV_X1 port map( A => ADD_WR(2), ZN => n14445);
   U16604 : INV_X1 port map( A => ADD_WR(0), ZN => n14447);
   U16605 : INV_X1 port map( A => ADD_WR(1), ZN => n14446);
   U16606 : INV_X1 port map( A => ADD_RD2(1), ZN => n14461);
   U16607 : INV_X1 port map( A => ADD_RD1(1), ZN => n14454);
   U16608 : INV_X1 port map( A => n16730, ZN => n16739);
   U16609 : INV_X1 port map( A => n16731, ZN => n16832);
   U16610 : CLKBUF_X1 port map( A => n14442, Z => n17320);

end SYN_A;
