
library IEEE;

use IEEE.std_logic_1164.all;

package 
   CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4 
   is

-- define attributes
attribute ENUM_ENCODING : STRING;

end 
   CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4.all;

entity control_unit is

   port( clock, reset, call, ret, mmu_ack : in std_logic;  cwp_out, swp_out : 
         out std_logic_vector (3 downto 0);  fill, spill : out std_logic);

end control_unit;

architecture SYN_Behavioral of control_unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal cwp_out_3_port, cwp_out_2_port, cwp_out_1_port, cwp_out_0_port, 
      swp_out_3_port, swp_out_2_port, swp_out_1_port, swp_out_0_port, N36, N39,
      cansave_3_port, cansave_2_port, cansave_1_port, cansave_0_port, 
      canrestore_3_port, canrestore_2_port, canrestore_1_port, 
      canrestore_0_port, N146, N148, N154, N156, N160, N162, N164, N166, N168, 
      N170, N172, N174, N176, N182, N186, N190, N198, N199, N28, 
      CurrState_2_port, CurrState_1_port, CurrState_0_port, n21, n24, n25, n26,
      n27, n36_port, n41, n57, n73, n76, n88, n63, n22, n23, n28_port, n29, n30
      , n31, n32, n33, n34, n35, n37, n38, n39_port, n40, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61
      , n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92 : 
      std_logic;

begin
   cwp_out <= ( cwp_out_3_port, cwp_out_2_port, cwp_out_1_port, cwp_out_0_port 
      );
   swp_out <= ( swp_out_3_port, swp_out_2_port, swp_out_1_port, swp_out_0_port 
      );
   
   canrestore_reg_0_inst : DLH_X1 port map( G => N198, D => N170, Q => 
                           canrestore_0_port);
   cansave_reg_3_inst : DLH_X1 port map( G => N198, D => N168, Q => 
                           cansave_3_port);
   fill_reg : DLH_X1 port map( G => N182, D => N39, Q => fill);
   cansave_reg_0_inst : DLH_X1 port map( G => N198, D => N162, Q => 
                           cansave_0_port);
   cansave_reg_1_inst : DLH_X1 port map( G => N198, D => N164, Q => 
                           cansave_1_port);
   cansave_reg_2_inst : DLH_X1 port map( G => N198, D => N166, Q => 
                           cansave_2_port);
   spill_reg : DLH_X1 port map( G => N199, D => N36, Q => spill);
   canrestore_reg_1_inst : DLH_X1 port map( G => N198, D => N172, Q => 
                           canrestore_1_port);
   canrestore_reg_2_inst : DLH_X1 port map( G => N198, D => N174, Q => 
                           canrestore_2_port);
   canrestore_reg_3_inst : DLH_X1 port map( G => N198, D => N176, Q => 
                           canrestore_3_port);
   cwp_reg_0_inst : DLH_X1 port map( G => N190, D => N154, Q => cwp_out_0_port)
                           ;
   swp_reg_0_inst : DLH_X1 port map( G => N186, D => N146, Q => swp_out_0_port)
                           ;
   swp_reg_1_inst : DLH_X1 port map( G => N186, D => N148, Q => swp_out_1_port)
                           ;
   cwp_reg_2_inst : DLH_X1 port map( G => N190, D => N160, Q => cwp_out_2_port)
                           ;
   cwp_reg_3_inst : DLH_X1 port map( G => N190, D => N160, Q => cwp_out_3_port)
                           ;
   cwp_reg_1_inst : DLH_X1 port map( G => N190, D => N156, Q => cwp_out_1_port)
                           ;
   U5 : AOI211_X2 port map( C1 => N36, C2 => n63, A => N39, B => n26, ZN => n21
                           );
   U6 : AND3_X2 port map( A1 => mmu_ack, A2 => N28, A3 => n27, ZN => n26);
   U25 : NAND2_X2 port map( A1 => n27, A2 => CurrState_0_port, ZN => n25);
   U26 : NOR2_X2 port map( A1 => n41, A2 => CurrState_1_port, ZN => n27);
   U38 : NOR3_X2 port map( A1 => CurrState_2_port, A2 => CurrState_0_port, A3 
                           => n57, ZN => N36);
   U87 : NOR2_X2 port map( A1 => n88, A2 => call, ZN => n76);
   U89 : NOR3_X2 port map( A1 => CurrState_2_port, A2 => CurrState_1_port, A3 
                           => N28, ZN => n36_port);
   U103 : NAND3_X1 port map( A1 => n41, A2 => n57, A3 => N28, ZN => n24);
   U106 : NAND3_X1 port map( A1 => CurrState_0_port, A2 => n41, A3 => 
                           CurrState_1_port, ZN => n73);
   swp_out_2_port <= '0';
   swp_out_3_port <= '0';
   U84 : XOR2_X1 port map( A => n38, B => n39_port, Z => n37);
   U85 : XOR2_X1 port map( A => canrestore_3_port, B => n40, Z => n39_port);
   U86 : XOR2_X1 port map( A => canrestore_2_port, B => n40, Z => n45);
   U88 : NAND3_X1 port map( A1 => n48, A2 => n51, A3 => canrestore_0_port, ZN 
                           => n50);
   U90 : XOR2_X1 port map( A => n54, B => n55, Z => n53);
   U91 : XOR2_X1 port map( A => cansave_3_port, B => n56, Z => n55);
   U92 : XOR2_X1 port map( A => n60, B => n64, Z => n62);
   U93 : XOR2_X1 port map( A => cansave_2_port, B => n56, Z => n64);
   U94 : NAND3_X1 port map( A1 => n66, A2 => n51, A3 => cansave_0_port, ZN => 
                           n68);
   U95 : XOR2_X1 port map( A => n56, B => cansave_1_port, Z => n66);
   U96 : NAND3_X1 port map( A1 => n70, A2 => n88, A3 => n73, ZN => n51);
   U97 : XOR2_X1 port map( A => swp_out_1_port, B => n23, Z => n77);
   U98 : NAND3_X1 port map( A1 => n28_port, A2 => n29, A3 => n27, ZN => n90);
   U3 : INV_X1 port map( A => n46, ZN => n40);
   U4 : NOR2_X1 port map( A1 => n52, A2 => n31, ZN => n46);
   U7 : INV_X1 port map( A => n61, ZN => n56);
   U8 : INV_X1 port map( A => n80, ZN => n75);
   U11 : OAI22_X1 port map( A1 => n78, A2 => n79, B1 => n80, B2 => n81, ZN => 
                           n74);
   U12 : NAND2_X1 port map( A1 => n84, A2 => n81, ZN => n78);
   U13 : INV_X1 port map( A => n85, ZN => n81);
   U14 : OAI22_X1 port map( A1 => n34, A2 => n23, B1 => n82, B2 => n83, ZN => 
                           n79);
   U15 : OAI22_X1 port map( A1 => n82, A2 => n83, B1 => n87, B2 => n89, ZN => 
                           n80);
   U16 : INV_X1 port map( A => n84, ZN => n87);
   U17 : NOR2_X1 port map( A1 => n34, A2 => n23, ZN => n89);
   U18 : OAI21_X1 port map( B1 => n86, B2 => n31, A => n28_port, ZN => n32);
   U19 : NOR2_X1 port map( A1 => n70, A2 => n63, ZN => n31);
   U20 : INV_X1 port map( A => n51, ZN => n35);
   U21 : INV_X1 port map( A => n86, ZN => n34);
   U22 : NAND2_X1 port map( A1 => n34, A2 => n69, ZN => n61);
   U23 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => N198);
   U24 : INV_X1 port map( A => N190, ZN => n33);
   U27 : INV_X1 port map( A => n57, ZN => CurrState_1_port);
   U28 : INV_X1 port map( A => n83, ZN => n52);
   U29 : INV_X1 port map( A => N28, ZN => CurrState_0_port);
   U30 : INV_X1 port map( A => CurrState_2_port, ZN => n41);
   U31 : INV_X1 port map( A => n58, ZN => n60);
   U32 : AND2_X1 port map( A1 => n42, A2 => n40, ZN => n43);
   U33 : NOR4_X1 port map( A1 => canrestore_3_port, A2 => n73, A3 => 
                           canrestore_2_port, A4 => n91, ZN => n86);
   U34 : OR2_X1 port map( A1 => canrestore_1_port, A2 => canrestore_0_port, ZN 
                           => n91);
   U35 : OAI211_X1 port map( C1 => ret, C2 => call, A => n36_port, B => 
                           n28_port, ZN => n57);
   U36 : OAI22_X1 port map( A1 => cansave_0_port, A2 => n61, B1 => 
                           cansave_1_port, B2 => n65, ZN => n58);
   U37 : AND2_X1 port map( A1 => n61, A2 => cansave_0_port, ZN => n65);
   U39 : OAI21_X1 port map( B1 => n46, B2 => n22, A => n47, ZN => n42);
   U40 : INV_X1 port map( A => canrestore_0_port, ZN => n22);
   U41 : OAI21_X1 port map( B1 => canrestore_0_port, B2 => n40, A => 
                           canrestore_1_port, ZN => n47);
   U42 : OAI21_X1 port map( B1 => reset, B2 => n24, A => n57, ZN => N190);
   U43 : OAI221_X1 port map( B1 => cwp_out_0_port, B2 => n69, C1 => n75, C2 => 
                           n72, A => n24, ZN => N154);
   U44 : OAI221_X1 port map( B1 => n71, B2 => n69, C1 => n72, C2 => n74, A => 
                           n24, ZN => N156);
   U45 : XNOR2_X1 port map( A => cwp_out_0_port, B => cwp_out_1_port, ZN => n71
                           );
   U46 : OAI22_X1 port map( A1 => swp_out_0_port, A2 => n70, B1 => n73, B2 => 
                           n75, ZN => N146);
   U47 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => n77, B2 => n70, ZN => 
                           N148);
   U48 : AOI22_X1 port map( A1 => n86, A2 => swp_out_1_port, B1 => 
                           cwp_out_1_port, B2 => n52, ZN => n85);
   U49 : NOR2_X1 port map( A1 => cwp_out_2_port, A2 => cwp_out_3_port, ZN => 
                           n82);
   U50 : NAND2_X1 port map( A1 => n28_port, A2 => n92, ZN => N28);
   U51 : NAND4_X1 port map( A1 => n25, A2 => n21, A3 => n24, A4 => n72, ZN => 
                           n92);
   U52 : NOR2_X1 port map( A1 => n35, A2 => canrestore_0_port, ZN => N170);
   U53 : NOR2_X1 port map( A1 => n35, A2 => cansave_0_port, ZN => N162);
   U54 : NAND2_X1 port map( A1 => n32, A2 => n90, ZN => CurrState_2_port);
   U55 : INV_X1 port map( A => mmu_ack, ZN => n29);
   U56 : OR4_X1 port map( A1 => cansave_0_port, A2 => cansave_1_port, A3 => 
                           cansave_2_port, A4 => cansave_3_port, ZN => n63);
   U57 : OAI21_X1 port map( B1 => n60, B2 => n61, A => cansave_2_port, ZN => 
                           n59);
   U58 : NAND2_X1 port map( A1 => ret, A2 => n76, ZN => n83);
   U59 : NAND2_X1 port map( A1 => call, A2 => n36_port, ZN => n69);
   U60 : INV_X1 port map( A => N36, ZN => n70);
   U61 : AOI21_X1 port map( B1 => n25, B2 => n34, A => reset, ZN => N182);
   U62 : INV_X1 port map( A => reset, ZN => n28_port);
   U63 : OAI21_X1 port map( B1 => reset, B2 => n24, A => n32, ZN => N186);
   U64 : INV_X1 port map( A => n73, ZN => N39);
   U65 : NAND2_X1 port map( A1 => n52, A2 => cwp_out_0_port, ZN => n84);
   U66 : INV_X1 port map( A => n76, ZN => n72);
   U67 : INV_X1 port map( A => swp_out_0_port, ZN => n23);
   U68 : INV_X1 port map( A => n36_port, ZN => n88);
   U69 : OAI21_X1 port map( B1 => n35, B2 => n62, A => n24, ZN => N166);
   U70 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => N164);
   U71 : INV_X1 port map( A => N162, ZN => n67);
   U72 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => N172);
   U73 : INV_X1 port map( A => N170, ZN => n49);
   U74 : XNOR2_X1 port map( A => canrestore_1_port, B => n40, ZN => n48);
   U75 : NOR2_X1 port map( A1 => n35, A2 => n37, ZN => N176);
   U76 : OAI22_X1 port map( A1 => n40, A2 => n42, B1 => canrestore_2_port, B2 
                           => n43, ZN => n38);
   U77 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => N174);
   U78 : XNOR2_X1 port map( A => n45, B => n42, ZN => n44);
   U79 : NOR2_X1 port map( A1 => n35, A2 => n53, ZN => N168);
   U80 : OAI21_X1 port map( B1 => n56, B2 => n58, A => n59, ZN => n54);
   U81 : NOR2_X1 port map( A1 => reset, A2 => n30, ZN => N199);
   U82 : AOI21_X1 port map( B1 => n27, B2 => N28, A => n31, ZN => n30);
   U83 : INV_X1 port map( A => n24, ZN => N160);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4.all;

entity register_file_NBIT32_NADDRESS5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT32_NADDRESS5;

architecture SYN_A of register_file_NBIT32_NADDRESS5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
      n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
      n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
      n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
      n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
      n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
      n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
      n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
      n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
      n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
      n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
      n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, 
      n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
      n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
      n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
      n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
      n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
      n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
      n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
      n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
      n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, 
      n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
      n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
      n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, 
      n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, 
      n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
      n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
      n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, 
      n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
      n2295, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
      n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
      n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
      n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, 
      n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
      n3255, n3256, n3257, n3258, n3259, n6315, n6316, n6317, n6318, n6319, 
      n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, 
      n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, 
      n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, 
      n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, 
      n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, 
      n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
      n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
      n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
      n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, 
      n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, 
      n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, 
      n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
      n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
      n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
      n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, 
      n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, 
      n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
      n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
      n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, 
      n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
      n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
      n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, 
      n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, 
      n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, 
      n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
      n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
      n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, 
      n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, 
      n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, 
      n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, 
      n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, 
      n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, 
      n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
      n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
      n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3263, n3264, n3265, 
      n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, 
      n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, 
      n3286, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3384, n3386, n3388, n3390, n3392, n3394, n3396, 
      n3398, n3400, n3402, n3404, n3406, n3408, n3410, n3412, n3414, n3416, 
      n3418, n3420, n3422, n3424, n3426, n3428, n3430, n3432, n3434, n3436, 
      n3438, n3440, n3442, n3444, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
      n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
      n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
      n3482, n3483, n3484, n3485, n3486, n3519, n3520, n3521, n3522, n3523, 
      n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, 
      n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, 
      n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
      n3554, n3555, n3556, n3557, n3558, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
      n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3599, 
      n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
      n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, 
      n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, 
      n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, 
      n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
      n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
      n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
      n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n7637, n7638, n7639, n7640, n7641, 
      n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, 
      n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
      n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, 
      n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, 
      n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, 
      n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, 
      n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, 
      n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, 
      n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, 
      n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, 
      n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, 
      n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, 
      n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, 
      n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, 
      n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, 
      n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, 
      n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
      n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, 
      n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, 
      n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, 
      n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, 
      n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, 
      n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, 
      n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, 
      n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, 
      n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, 
      n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, 
      n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, 
      n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, 
      n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, 
      n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, 
      n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, 
      n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, 
      n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, 
      n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, 
      n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, 
      n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, 
      n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, 
      n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, 
      n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, 
      n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, 
      n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, 
      n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, 
      n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, 
      n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, 
      n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, 
      n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, 
      n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, 
      n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, 
      n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, 
      n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, 
      n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, 
      n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, 
      n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, 
      n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, 
      n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, 
      n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, 
      n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, 
      n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, 
      n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, 
      n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, 
      n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, 
      n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, 
      n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, 
      n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, 
      n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, 
      n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, 
      n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, 
      n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, 
      n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, 
      n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, 
      n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, 
      n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, 
      n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, 
      n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, 
      n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, 
      n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, 
      n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, 
      n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, 
      n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, 
      n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, 
      n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, 
      n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, 
      n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, 
      n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, 
      n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, 
      n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, 
      n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, 
      n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, 
      n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, 
      n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, 
      n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, 
      n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, 
      n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, 
      n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, 
      n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, 
      n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, 
      n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, 
      n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, 
      n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, 
      n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, 
      n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, 
      n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, 
      n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, 
      n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, 
      n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, 
      n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, 
      n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, 
      n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, 
      n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, 
      n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, 
      n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, 
      n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, 
      n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, 
      n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, 
      n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, 
      n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, 
      n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, 
      n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, 
      n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, 
      n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, 
      n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, 
      n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, 
      n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, 
      n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, 
      n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, 
      n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, 
      n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, 
      n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, 
      n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, 
      n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, 
      n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, 
      n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, 
      n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, 
      n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, 
      n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, 
      n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, 
      n9022, n9023, n9024, n9025, n_1000, n_1001, n_1002, n_1003, n_1004, 
      n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, 
      n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => n3622
                           , QN => n7916);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => n3621
                           , QN => n7915);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => n3620
                           , QN => n7914);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => n3619
                           , QN => n7913);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => n3618
                           , QN => n7912);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => n3617
                           , QN => n7911);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => n3616
                           , QN => n7910);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => n3615
                           , QN => n7909);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => n3862
                           , QN => n8204);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => n3861
                           , QN => n8203);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => n3860
                           , QN => n8202);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => n3859
                           , QN => n8201);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => n3858
                           , QN => n8200);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => n3857
                           , QN => n8199);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => n3856
                           , QN => n8198);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => n3855
                           , QN => n8197);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => n3854
                           , QN => n8196);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => n3853
                           , QN => n8195);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => n3852
                           , QN => n8194);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => n3851
                           , QN => n8193);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => n3850
                           , QN => n8192);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => n3849
                           , QN => n8191);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => n3848,
                           QN => n8190);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => n3847,
                           QN => n8189);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => n3846,
                           QN => n8188);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => n3845,
                           QN => n8187);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => n3844,
                           QN => n8186);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => n3843,
                           QN => n8185);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => n3842,
                           QN => n8184);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => n3841,
                           QN => n8183);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => n3840,
                           QN => n8182);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => n3839,
                           QN => n8181);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => n3614
                           , QN => n7868);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => n3613
                           , QN => n7867);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => n3612
                           , QN => n7866);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => n3611
                           , QN => n7865);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => n3610
                           , QN => n7864);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => n3609
                           , QN => n7863);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => n3608
                           , QN => n7862);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => n3607
                           , QN => n7861);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => n3838
                           , QN => n8132);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => n3837
                           , QN => n8131);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => n3836
                           , QN => n8130);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => n3835
                           , QN => n8129);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => n3834
                           , QN => n8128);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => n3833
                           , QN => n8127);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => n3832
                           , QN => n8126);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => n3831
                           , QN => n8125);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => n3830
                           , QN => n8124);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => n3829
                           , QN => n8123);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => n3828
                           , QN => n8122);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => n3827
                           , QN => n8121);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => n3826
                           , QN => n8120);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => n3825
                           , QN => n8119);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => n3824,
                           QN => n8118);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => n3823,
                           QN => n8117);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => n3822,
                           QN => n8116);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => n3821,
                           QN => n8115);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => n3820,
                           QN => n8114);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => n3819,
                           QN => n8113);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => n3818,
                           QN => n8112);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => n3817,
                           QN => n8111);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => n3816,
                           QN => n8110);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => n3815,
                           QN => n8109);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => n6602
                           , QN => n7644);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => n6601
                           , QN => n7643);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => n6600
                           , QN => n7642);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => n6599
                           , QN => n7641);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => n6598
                           , QN => n7640);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => n6597
                           , QN => n7639);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => n6596
                           , QN => n7638);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => n6595
                           , QN => n7637);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => n6594
                           , QN => n7656);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => n6593
                           , QN => n7655);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => n6592
                           , QN => n7654);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => n6591
                           , QN => n7653);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => n6590
                           , QN => n7652);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => n6589
                           , QN => n7651);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => n6588
                           , QN => n7650);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => n6587
                           , QN => n7649);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => n6586
                           , QN => n7648);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => n6585
                           , QN => n7647);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => n6584
                           , QN => n7646);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => n6583
                           , QN => n7645);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => n6582
                           , QN => n7740);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => n6581
                           , QN => n7739);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => n6580,
                           QN => n7738);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => n6579,
                           QN => n7737);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => n6578,
                           QN => n7736);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => n6577,
                           QN => n7735);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => n6576,
                           QN => n7734);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => n6575,
                           QN => n7733);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => n6574,
                           QN => n7732);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => n6573,
                           QN => n7731);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => n6572,
                           QN => n7730);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => n6571,
                           QN => n7729);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => n3606
                           , QN => n7760);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => n3605
                           , QN => n7759);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => n3604
                           , QN => n7758);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => n3603
                           , QN => n7757);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => n3602
                           , QN => n7756);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => n3601
                           , QN => n7755);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => n3600
                           , QN => n7754);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => n3599
                           , QN => n7753);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => n3814
                           , QN => n7752);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => n3813
                           , QN => n7751);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => n3812
                           , QN => n7750);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => n3811
                           , QN => n7749);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => n3810
                           , QN => n7748);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => n3809
                           , QN => n7747);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => n3808
                           , QN => n7746);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => n3807
                           , QN => n7745);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => n3806
                           , QN => n7744);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => n3805
                           , QN => n7743);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => n3804
                           , QN => n7742);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => n3803
                           , QN => n7741);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => n3802
                           , QN => n7888);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => n3801
                           , QN => n7887);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => n3800,
                           QN => n7886);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n3799,
                           QN => n7885);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => n3798,
                           QN => n7884);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => n3797,
                           QN => n7883);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => n3796,
                           QN => n7882);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => n3795,
                           QN => n7881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => n3794,
                           QN => n7880);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => n3793,
                           QN => n7879);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => n3792,
                           QN => n7878);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => n3791,
                           QN => n7877);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => n3286
                           , QN => n7972);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => n3285
                           , QN => n7971);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => n3284
                           , QN => n7970);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => n3283
                           , QN => n7969);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => n3282
                           , QN => n7968);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => n3281
                           , QN => n7967);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => n3280
                           , QN => n7966);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => n3279
                           , QN => n7965);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => n3382
                           , QN => n8436);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => n3381
                           , QN => n8435);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => n3380
                           , QN => n8434);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => n3379
                           , QN => n8433);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => n3378
                           , QN => n8432);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => n3377
                           , QN => n8431);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => n3376
                           , QN => n8430);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => n3375
                           , QN => n8429);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => n3374
                           , QN => n8428);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => n3373
                           , QN => n8427);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => n3372
                           , QN => n8426);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => n3371
                           , QN => n8425);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => n3370
                           , QN => n8424);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => n3369
                           , QN => n8423);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => n3368,
                           QN => n8422);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n3367,
                           QN => n8421);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => n3366,
                           QN => n8420);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => n3365,
                           QN => n8419);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => n3364,
                           QN => n8418);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => n3363,
                           QN => n8417);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => n3362,
                           QN => n8416);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => n3361,
                           QN => n8415);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => n3360,
                           QN => n8414);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => n3359,
                           QN => n8413);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => n8260
                           , QN => n6810);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => n8259
                           , QN => n6809);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => n8258
                           , QN => n6808);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => n8257
                           , QN => n6807);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => n8256
                           , QN => n6806);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => n8255
                           , QN => n6805);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => n8254
                           , QN => n6804);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => n8253
                           , QN => n6803);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => n8252
                           , QN => n6858);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => n8251
                           , QN => n6857);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => n8250
                           , QN => n6856);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => n8249
                           , QN => n6855);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => n8248
                           , QN => n6854);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => n8247
                           , QN => n6853);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => n8246
                           , QN => n6852);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => n8245
                           , QN => n6851);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => n8244
                           , QN => n6850);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => n8243
                           , QN => n6849);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => n8242
                           , QN => n6848);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => n8241
                           , QN => n6847);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => n8240
                           , QN => n6846);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => n8239
                           , QN => n6845);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => n8238,
                           QN => n6844);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n8237,
                           QN => n6843);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => n8236,
                           QN => n6842);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => n8235,
                           QN => n6841);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => n8234,
                           QN => n6840);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => n8233,
                           QN => n6839);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => n8232,
                           QN => n6838);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => n8231,
                           QN => n6837);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => n8230,
                           QN => n6836);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => n8229,
                           QN => n6835);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => n3278
                           , QN => n7876);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => n3277
                           , QN => n7875);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => n3276
                           , QN => n7874);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => n3275
                           , QN => n7873);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => n3274
                           , QN => n7872);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => n3273
                           , QN => n7871);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => n3272
                           , QN => n7870);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => n3271
                           , QN => n7869);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => n3358
                           , QN => n8156);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => n3357
                           , QN => n8155);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => n3356
                           , QN => n8154);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => n3355
                           , QN => n8153);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => n3354
                           , QN => n8152);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => n3353
                           , QN => n8151);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => n3352
                           , QN => n8150);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => n3351
                           , QN => n8149);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => n3350
                           , QN => n8148);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => n3349
                           , QN => n8147);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => n3348
                           , QN => n8146);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => n3347
                           , QN => n8145);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => n3346
                           , QN => n8144);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => n3345
                           , QN => n8143);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => n3344,
                           QN => n8142);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n3343,
                           QN => n8141);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n3342,
                           QN => n8140);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n3341,
                           QN => n8139);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => n3340,
                           QN => n8138);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => n3339,
                           QN => n8137);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => n3338,
                           QN => n8136);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => n3337,
                           QN => n8135);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => n3336,
                           QN => n8134);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => n3335,
                           QN => n8133);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           n_1000, QN => n7820);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n_1001, QN => n7818);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n_1002, QN => n7816);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           n_1003, QN => n7814);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           n_1004, QN => n7812);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           n_1005, QN => n7810);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           n_1006, QN => n7808);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           n_1007, QN => n7806);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           n_1008, QN => n7679);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           n_1009, QN => n7677);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           n_1010, QN => n7675);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           n_1011, QN => n7673);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           n_1012, QN => n7671);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           n_1013, QN => n7669);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           n_1014, QN => n7667);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           n_1015, QN => n7665);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           n_1016, QN => n7663);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           n_1017, QN => n7661);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           n_1018, QN => n7659);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           n_1019, QN => n7657);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           n_1020, QN => n7803);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           n_1021, QN => n7801);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => n_1022
                           , QN => n7799);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n_1023
                           , QN => n7797);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => n_1024
                           , QN => n7796);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => n_1025
                           , QN => n7795);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => n_1026
                           , QN => n7794);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => n_1027
                           , QN => n7793);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => n_1028
                           , QN => n7792);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => n_1029
                           , QN => n7791);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => n_1030
                           , QN => n7790);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => n_1031
                           , QN => n7789);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => n3590
                           , QN => n7704);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => n3589
                           , QN => n7703);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => n3588
                           , QN => n7702);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => n3587
                           , QN => n7701);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => n3586
                           , QN => n7700);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => n3585
                           , QN => n7699);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => n3584
                           , QN => n7698);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => n3583
                           , QN => n7697);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => n3694
                           , QN => n7728);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => n3693
                           , QN => n7727);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => n3692
                           , QN => n7726);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => n3691
                           , QN => n7725);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => n3690
                           , QN => n7724);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => n3689
                           , QN => n7723);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => n3688
                           , QN => n7722);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => n3687
                           , QN => n7721);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => n3686
                           , QN => n7720);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => n3685
                           , QN => n7719);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => n3684
                           , QN => n7718);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => n3683
                           , QN => n7717);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => n3682
                           , QN => n7852);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => n3681
                           , QN => n7851);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => n3680,
                           QN => n7850);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => n3679,
                           QN => n7849);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => n3678,
                           QN => n7848);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => n3677,
                           QN => n7847);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => n3676,
                           QN => n7846);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => n3675,
                           QN => n7845);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => n3674,
                           QN => n7844);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => n3673,
                           QN => n7843);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => n3672,
                           QN => n7842);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => n3671,
                           QN => n7841);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           n_1032, QN => n6874);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n_1033, QN => n6873);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n_1034, QN => n6872);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n_1035, QN => n6871);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n_1036, QN => n6870);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n_1037, QN => n6869);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n_1038, QN => n6868);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n_1039, QN => n6867);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n_1040, QN => n6922);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n_1041, QN => n6921);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n_1042, QN => n6920);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n_1043, QN => n6919);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n_1044, QN => n6918);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n_1045, QN => n6917);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n_1046, QN => n6916);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n_1047, QN => n6915);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n_1048, QN => n6914);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n_1049, QN => n6913);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n_1050, QN => n6912);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n_1051, QN => n6911);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n_1052, QN => n6910);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n_1053, QN => n6909);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => n_1054
                           , QN => n6908);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => n_1055
                           , QN => n6907);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => n_1056
                           , QN => n6906);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => n_1057
                           , QN => n6905);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => n_1058
                           , QN => n6904);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => n_1059
                           , QN => n6903);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => n_1060
                           , QN => n6902);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => n_1061
                           , QN => n6901);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => n_1062
                           , QN => n6900);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => n_1063
                           , QN => n6899);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n3582, QN => n7768);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n3581, QN => n7767);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n3580, QN => n7766);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n3579, QN => n7765);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n3578, QN => n7764);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n3577, QN => n7763);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n3576, QN => n7762);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n3575, QN => n7761);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n3670, QN => n7780);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n3669, QN => n7779);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n3668, QN => n7778);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n3667, QN => n7777);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n3666, QN => n7776);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n3665, QN => n7775);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           n3664, QN => n7774);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           n3663, QN => n7773);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           n3662, QN => n7772);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           n3661, QN => n7771);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           n3660, QN => n7770);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           n3659, QN => n7769);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           n3658, QN => n7900);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           n3657, QN => n7899);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => n3656
                           , QN => n7898);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => n3655
                           , QN => n7897);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => n3654
                           , QN => n7896);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => n3653
                           , QN => n7895);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => n3652
                           , QN => n7894);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => n3651
                           , QN => n7893);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => n3650
                           , QN => n7892);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => n3649
                           , QN => n7891);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => n3648
                           , QN => n7890);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => n3647
                           , QN => n7889);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n3574, QN => n7964);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n3573, QN => n7963);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n3572, QN => n7962);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           n3571, QN => n7961);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           n3570, QN => n7960);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           n3569, QN => n7959);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           n3568, QN => n7958);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           n3567, QN => n7957);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           n3790, QN => n8412);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           n3789, QN => n8411);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           n3788, QN => n8410);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           n3787, QN => n8409);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           n3786, QN => n8408);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n3785, QN => n8407);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           n3784, QN => n8406);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           n3783, QN => n8405);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           n3782, QN => n8404);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           n3781, QN => n8403);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           n3780, QN => n8402);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           n3779, QN => n8401);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           n3778, QN => n8400);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           n3777, QN => n8399);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => n3776
                           , QN => n8398);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => n3775
                           , QN => n8397);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => n3774
                           , QN => n8396);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => n3773
                           , QN => n8395);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => n3772
                           , QN => n8394);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => n3771
                           , QN => n8393);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => n3770
                           , QN => n8392);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => n3769
                           , QN => n8391);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => n3768
                           , QN => n8390);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => n3767
                           , QN => n8389);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n8292, QN => n6746);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n8291, QN => n6745);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n8290, QN => n6744);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n8289, QN => n6743);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n8288, QN => n6742);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n8287, QN => n6741);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n8286, QN => n6740);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n8285, QN => n6739);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n8284, QN => n6794);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n8283, QN => n6793);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n8282, QN => n6792);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n8281, QN => n6791);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n8280, QN => n6790);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n8279, QN => n6789);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n8278, QN => n6788);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n8277, QN => n6787);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n8276, QN => n6786);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n8275, QN => n6785);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n8274, QN => n6784);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n8273, QN => n6783);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n8272, QN => n6782);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n8271, QN => n6781);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => n8270
                           , QN => n6780);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => n8269
                           , QN => n6779);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => n8268
                           , QN => n6778);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => n8267
                           , QN => n6777);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => n8266
                           , QN => n6776);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => n8265
                           , QN => n6775);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => n8264
                           , QN => n6774);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => n8263
                           , QN => n6773);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => n8262
                           , QN => n6772);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => n8261
                           , QN => n6771);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n_1064, QN => n6738);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n_1065, QN => n6737);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n_1066, QN => n6736);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n_1067, QN => n6735);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n_1068, QN => n6734);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n_1069, QN => n6733);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n_1070, QN => n6732);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n_1071, QN => n6731);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n_1072, QN => n6770);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n_1073, QN => n6769);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n_1074, QN => n6768);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n_1075, QN => n6767);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n_1076, QN => n6766);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n_1077, QN => n6765);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n_1078, QN => n6764);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n_1079, QN => n6763);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n_1080, QN => n6762);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n_1081, QN => n6761);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n_1082, QN => n6760);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n_1083, QN => n6759);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n_1084, QN => n6758);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n_1085, QN => n6757);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n_1086, QN => n6756);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n_1087, QN => n6755);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n_1088, QN => n6754);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n_1089, QN => n6753);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n_1090, QN => n6752);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n_1091, QN => n6751);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n_1092, QN => n6750);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n_1093, QN => n6749);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n_1094, QN => n6748);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n_1095, QN => n6747);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n8084, QN => n6802);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n8083, QN => n6801);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n8082, QN => n6800);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n8081, QN => n6799);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n8080, QN => n6798);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n8079, QN => n6797);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n8078, QN => n6796);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n8077, QN => n6795);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n8076, QN => n6834);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n8075, QN => n6833);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n8074, QN => n6832);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n8073, QN => n6831);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n8072, QN => n6830);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n8071, QN => n6829);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n8070, QN => n6828);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n8069, QN => n6827);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n8068, QN => n6826);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n8067, QN => n6825);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           n8066, QN => n6824);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           n8065, QN => n6823);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           n8064, QN => n6822);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           n8063, QN => n6821);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => n8062
                           , QN => n6820);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => n8061
                           , QN => n6819);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => n8060
                           , QN => n6818);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => n8059
                           , QN => n6817);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => n8058
                           , QN => n6816);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => n8057
                           , QN => n6815);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => n8056
                           , QN => n6814);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => n8055
                           , QN => n6813);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => n8054
                           , QN => n6812);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => n8053
                           , QN => n6811);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n_1096, QN => n7688);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n_1097, QN => n7687);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n_1098, QN => n7686);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n_1099, QN => n7685);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n_1100, QN => n7684);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n_1101, QN => n7683);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n_1102, QN => n7682);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n_1103, QN => n7681);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n_1104, QN => n7680);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n_1105, QN => n7678);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n_1106, QN => n7676);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n_1107, QN => n7674);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n_1108, QN => n7672);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n_1109, QN => n7670);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n_1110, QN => n7668);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n_1111, QN => n7666);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n_1112, QN => n7664);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n_1113, QN => n7662);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n_1114, QN => n7660);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n_1115, QN => n7658);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n_1116, QN => n7804);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n_1117, QN => n7802);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n_1118, QN => n7800);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           n_1119, QN => n7798);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           n_1120, QN => n7788);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           n_1121, QN => n7787);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           n_1122, QN => n7786);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           n_1123, QN => n7785);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n_1124, QN => n7784);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n_1125, QN => n7783);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n_1126, QN => n7782);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n_1127, QN => n7781);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n3558, QN => n7696);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n3557, QN => n7695);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n3556, QN => n7694);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n3555, QN => n7693);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n3554, QN => n7692);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n3553, QN => n7691);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n3552, QN => n7690);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n3551, QN => n7689);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n3646, QN => n7716);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n3645, QN => n7715);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n3644, QN => n7714);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n3643, QN => n7713);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n3642, QN => n7712);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n3641, QN => n7711);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n3640, QN => n7710);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n3639, QN => n7709);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n3638, QN => n7708);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n3637, QN => n7707);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           n3636, QN => n7706);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           n3635, QN => n7705);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           n3634, QN => n7840);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           n3633, QN => n7839);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => n3632
                           , QN => n7838);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => n3631
                           , QN => n7837);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => n3630
                           , QN => n7836);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => n3629
                           , QN => n7835);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => n3628
                           , QN => n7834);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => n3627
                           , QN => n7833);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => n3626
                           , QN => n7832);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => n3625
                           , QN => n7831);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => n3624
                           , QN => n7830);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => n3623
                           , QN => n7829);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n3550, QN => n7860);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n3549, QN => n7859);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n3548, QN => n7858);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n3547, QN => n7857);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n3546, QN => n7856);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n3545, QN => n7855);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n3544, QN => n7854);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n3543, QN => n7853);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n3742, QN => n8108);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n3741, QN => n8107);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n3740, QN => n8106);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n3739, QN => n8105);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n3738, QN => n8104);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n3737, QN => n8103);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n3736, QN => n8102);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n3735, QN => n8101);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n3734, QN => n8100);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n3733, QN => n8099);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n3732, QN => n8098);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n3731, QN => n8097);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n3730, QN => n8096);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n3729, QN => n8095);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => n3728
                           , QN => n8094);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => n3727
                           , QN => n8093);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => n3726
                           , QN => n8092);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => n3725
                           , QN => n8091);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => n3724
                           , QN => n8090);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => n3723
                           , QN => n8089);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => n3722
                           , QN => n8088);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => n3721
                           , QN => n8087);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => n3720
                           , QN => n8086);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => n3719
                           , QN => n8085);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n_1128, QN => n6682);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1129, QN => n6681);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1130, QN => n6680);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1131, QN => n6679);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1132, QN => n6678);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1133, QN => n6677);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1134, QN => n6676);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1135, QN => n6675);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1136, QN => n6730);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1137, QN => n6729);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1138, QN => n6728);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1139, QN => n6727);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1140, QN => n6726);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1141, QN => n6725);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1142, QN => n6724);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1143, QN => n6723);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1144, QN => n6722);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1145, QN => n6721);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1146, QN => n6720);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1147, QN => n6719);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1148, QN => n6718);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1149, QN => n6717);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1150, QN => n6716);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1151, QN => n6715);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n_1152, QN => n6714);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n_1153, QN => n6713);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n_1154, QN => n6712);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n_1155, QN => n6711);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1156, QN => n6710);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1157, QN => n6709);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1158, QN => n6708);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1159, QN => n6707);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n3542, QN => n7940);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n3541, QN => n7939);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n3540, QN => n7938);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n3539, QN => n7937);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n3538, QN => n7936);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n3537, QN => n7935);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n3536, QN => n7934);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n3535, QN => n7933);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n3534, QN => n8340);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n3533, QN => n8339);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n3532, QN => n8338);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n3531, QN => n8337);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n3530, QN => n8336);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n3529, QN => n8335);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n3528, QN => n8334);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n3527, QN => n8333);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n3526, QN => n8332);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n3525, QN => n8331);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n3524, QN => n8330);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n3523, QN => n8329);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n3522, QN => n8328);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n3521, QN => n8327);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => n3520
                           , QN => n8326);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => n3519
                           , QN => n8325);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => n3486
                           , QN => n8324);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => n3485
                           , QN => n8323);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => n3484
                           , QN => n8322);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => n3483
                           , QN => n8321);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => n3482
                           , QN => n8320);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => n3481
                           , QN => n8319);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => n3480
                           , QN => n8318);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => n3479
                           , QN => n8317);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n3270, QN => n7924);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n3269, QN => n7923);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n3268, QN => n7922);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n3267, QN => n7921);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n3266, QN => n7920);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n3265, QN => n7919);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n3264, QN => n7918);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n3263, QN => n7917);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n3334, QN => n8228);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n3333, QN => n8227);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n3332, QN => n8226);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n3331, QN => n8225);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n3330, QN => n8224);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n3329, QN => n8223);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n3328, QN => n8222);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n3327, QN => n8221);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n3326, QN => n8220);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n3325, QN => n8219);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n3324, QN => n8218);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n3323, QN => n8217);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n3322, QN => n8216);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n3321, QN => n8215);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => n3320
                           , QN => n8214);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => n3319
                           , QN => n8213);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => n3318
                           , QN => n8212);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => n3317
                           , QN => n8211);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => n3316
                           , QN => n8210);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n3315
                           , QN => n8209);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => n3314
                           , QN => n8208);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n3313
                           , QN => n8207);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => n3312
                           , QN => n8206);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n3311
                           , QN => n8205);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n_1160, QN => n6338);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n_1161, QN => n6337);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n_1162, QN => n6336);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n_1163, QN => n6335);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n_1164, QN => n6334);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n_1165, QN => n6333);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n_1166, QN => n6332);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n_1167, QN => n6331);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n_1168, QN => n6330);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n_1169, QN => n6329);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n_1170, QN => n6328);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n_1171, QN => n6327);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n_1172, QN => n6326);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n_1173, QN => n6325);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n_1174, QN => n6324);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n_1175, QN => n6323);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n_1176, QN => n6322);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n_1177, QN => n6321);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n_1178, QN => n6320);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n_1179, QN => n6319);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n_1180, QN => n6318);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n_1181, QN => n6317);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n_1182, QN => n6316);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           n_1183, QN => n6315);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n_1184, QN => n6346);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           n_1185, QN => n6345);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n_1186, QN => n6344);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           n_1187, QN => n6343);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n_1188, QN => n6342);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           n_1189, QN => n6341);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n_1190, QN => n6340);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           n_1191, QN => n6339);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n_1192, QN => n7819);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n_1193, QN => n7817);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n_1194, QN => n7815);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n_1195, QN => n7813);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n_1196, QN => n7811);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n_1197, QN => n7809);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n_1198, QN => n7807);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n_1199, QN => n7805);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n_1200, QN => n7996);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n_1201, QN => n7995);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n_1202, QN => n7994);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n_1203, QN => n7993);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n_1204, QN => n7992);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n_1205, QN => n7991);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n_1206, QN => n7990);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n_1207, QN => n7989);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n_1208, QN => n7988);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n_1209, QN => n7987);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n_1210, QN => n7986);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n_1211, QN => n7985);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n_1212, QN => n7984);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n_1213, QN => n7983);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n_1214, QN => n7982);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           n_1215, QN => n7981);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n_1216, QN => n7980);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           n_1217, QN => n7979);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n_1218, QN => n7978);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           n_1219, QN => n7977);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n_1220, QN => n7976);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           n_1221, QN => n7975);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n_1222, QN => n7974);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           n_1223, QN => n7973);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n3446, QN => n7932);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n3444, QN => n7931);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n3442, QN => n7930);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n3440, QN => n7929);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n3438, QN => n7928);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n3436, QN => n7927);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n3434, QN => n7926);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n3432, QN => n7925);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n3430, QN => n8316);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n3428, QN => n8315);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n3426, QN => n8314);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n3424, QN => n8313);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n3422, QN => n8312);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n3420, QN => n8311);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n3418, QN => n8310);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n3416, QN => n8309);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n3414, QN => n8308);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n3412, QN => n8307);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n3410, QN => n8306);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n3408, QN => n8305);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n3406, QN => n8304);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n3404, QN => n8303);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => n3402
                           , QN => n8302);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n3400
                           , QN => n8301);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => n3398
                           , QN => n8300);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n3396
                           , QN => n8299);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => n3394
                           , QN => n8298);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n3392
                           , QN => n8297);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => n3390
                           , QN => n8296);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n3388
                           , QN => n8295);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => n3386
                           , QN => n8294);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n3384
                           , QN => n8293);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n_1224, QN => n6866);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n_1225, QN => n6865);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n_1226, QN => n6864);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n_1227, QN => n6863);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n_1228, QN => n6862);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n_1229, QN => n6861);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n_1230, QN => n6860);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n_1231, QN => n6859);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n_1232, QN => n6898);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n_1233, QN => n6897);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n_1234, QN => n6896);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n_1235, QN => n6895);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n_1236, QN => n6894);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n_1237, QN => n6893);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n_1238, QN => n6892);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n_1239, QN => n6891);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n_1240, QN => n6890);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n_1241, QN => n6889);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n_1242, QN => n6888);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n_1243, QN => n6887);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n_1244, QN => n6886);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n_1245, QN => n6885);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n_1246, QN => n6884);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n_1247, QN => n6883);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n_1248, QN => n6882);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n_1249, QN => n6881);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n_1250, QN => n6880);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n_1251, QN => n6879);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n_1252, QN => n6878);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n_1253, QN => n6877);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n_1254, QN => n6876);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n_1255, QN => n6875);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n3478, QN => n7908);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n3477, QN => n7907);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n3476, QN => n7906);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n3475, QN => n7905);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n3474, QN => n7904);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n3473, QN => n7903);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n3472, QN => n7902);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n3471, QN => n7901);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n3470, QN => n8180);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n3469, QN => n8179);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n3468, QN => n8178);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n3467, QN => n8177);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n3466, QN => n8176);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n3465, QN => n8175);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           n3464, QN => n8174);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           n3463, QN => n8173);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           n3462, QN => n8172);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           n3461, QN => n8171);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           n3460, QN => n8170);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           n3459, QN => n8169);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           n3458, QN => n8168);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           n3457, QN => n8167);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n3456
                           , QN => n8166);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n3455
                           , QN => n8165);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n3454
                           , QN => n8164);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n3453
                           , QN => n8163);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n3452
                           , QN => n8162);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n3451
                           , QN => n8161);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n3450
                           , QN => n8160);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n3449
                           , QN => n8159);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n3448
                           , QN => n8158);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n3447
                           , QN => n8157);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n_1256, QN => n6674);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n_1257, QN => n6673);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n_1258, QN => n6672);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n_1259, QN => n6671);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n_1260, QN => n6670);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n_1261, QN => n6669);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n_1262, QN => n6668);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n_1263, QN => n6667);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n_1264, QN => n6706);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n_1265, QN => n6705);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n_1266, QN => n6704);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n_1267, QN => n6703);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n_1268, QN => n6702);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n_1269, QN => n6701);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n_1270, QN => n6700);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n_1271, QN => n6699);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n_1272, QN => n6698);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n_1273, QN => n6697);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n_1274, QN => n6696);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n_1275, QN => n6695);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n_1276, QN => n6694);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n_1277, QN => n6693);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n_1278, QN => n6692);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n_1279, QN => n6691);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n_1280, QN => n6690);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n_1281, QN => n6689);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n_1282, QN => n6688);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n_1283, QN => n6687);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n_1284, QN => n6686);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n_1285, QN => n6685);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n_1286, QN => n6684);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n_1287, QN => n6683);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n_1288, QN => n7828);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n_1289, QN => n7827);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n_1290, QN => n7826);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n_1291, QN => n7825);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n_1292, QN => n7824);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n_1293, QN => n7823);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n_1294, QN => n7822);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n_1295, QN => n7821);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n_1296, QN => n8052);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n_1297, QN => n8051);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n_1298, QN => n8050);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n_1299, QN => n8049);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n_1300, QN => n8048);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n_1301, QN => n8047);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n_1302, QN => n8046);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n_1303, QN => n8045);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n_1304, QN => n8044);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n_1305, QN => n8043);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n_1306, QN => n8042);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n_1307, QN => n8041);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n_1308, QN => n8040);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n_1309, QN => n8039);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n_1310, QN => n8038);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n_1311, QN => n8037);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n_1312, QN => n8036);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n_1313, QN => n8035);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n_1314, QN => n8034);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n_1315, QN => n8033);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n_1316, QN => n8032);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n_1317, QN => n8031);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n_1318, QN => n8030);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n_1319, QN => n8029);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n6378, QN => n7956);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n6377, QN => n7955);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n6376, QN => n7954);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n6375, QN => n7953);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n6374, QN => n7952);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n6373, QN => n7951);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n6372, QN => n7950);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n6371, QN => n7949);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n6370, QN => n8388);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n6369, QN => n8387);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n6368, QN => n8386);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n6367, QN => n8385);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n6366, QN => n8384);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n6365, QN => n8383);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           n6364, QN => n8382);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           n6363, QN => n8381);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           n6362, QN => n8380);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           n6361, QN => n8379);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           n6360, QN => n8378);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           n6359, QN => n8377);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           n6358, QN => n8376);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           n6357, QN => n8375);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n6356
                           , QN => n8374);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n6355
                           , QN => n8373);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n6354
                           , QN => n8372);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n6353
                           , QN => n8371);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n6352
                           , QN => n8370);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n6351
                           , QN => n8369);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n6350
                           , QN => n8368);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n6349
                           , QN => n8367);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n6348
                           , QN => n8366);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n6347
                           , QN => n8365);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           n6666, QN => n7948);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n6665, QN => n7947);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n6664, QN => n7946);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n6663, QN => n7945);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n6662, QN => n7944);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n6661, QN => n7943);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n6660, QN => n7942);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n6659, QN => n7941);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n6658, QN => n8364);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n6657, QN => n8363);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n6656, QN => n8362);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n6655, QN => n8361);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n6654, QN => n8360);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n6653, QN => n8359);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           n6652, QN => n8358);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           n6651, QN => n8357);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           n6650, QN => n8356);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           n6649, QN => n8355);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           n6648, QN => n8354);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           n6647, QN => n8353);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           n6646, QN => n8352);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           n6645, QN => n8351);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n6644
                           , QN => n8350);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n6643
                           , QN => n8349);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n6642
                           , QN => n8348);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n6641
                           , QN => n8347);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n6640
                           , QN => n8346);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n6639
                           , QN => n8345);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n6638
                           , QN => n8344);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n6637
                           , QN => n8343);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n6636
                           , QN => n8342);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n6635
                           , QN => n8341);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           n_1320, QN => n6626);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           n_1321, QN => n6625);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           n_1322, QN => n6624);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           n_1323, QN => n6623);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           n_1324, QN => n6622);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           n_1325, QN => n6621);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           n_1326, QN => n6620);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           n_1327, QN => n6619);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           n_1328, QN => n6618);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           n_1329, QN => n6617);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           n_1330, QN => n6616);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           n_1331, QN => n6615);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           n_1332, QN => n6614);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           n_1333, QN => n6613);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           n_1334, QN => n6612);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           n_1335, QN => n6611);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           n_1336, QN => n6610);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           n_1337, QN => n6609);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           n_1338, QN => n6608);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           n_1339, QN => n6607);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           n_1340, QN => n6606);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           n_1341, QN => n6605);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           n_1342, QN => n6604);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           n_1343, QN => n6603);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           n_1344, QN => n6634);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           n_1345, QN => n6633);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           n_1346, QN => n6632);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           n_1347, QN => n6631);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           n_1348, QN => n6630);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           n_1349, QN => n6629);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           n_1350, QN => n6628);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           n_1351, QN => n6627);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           n_1352, QN => n8028);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           n_1353, QN => n8027);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           n_1354, QN => n8026);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           n_1355, QN => n8025);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           n_1356, QN => n8024);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           n_1357, QN => n8023);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           n_1358, QN => n8022);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           n_1359, QN => n8021);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           n_1360, QN => n8020);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           n_1361, QN => n8019);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           n_1362, QN => n8018);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           n_1363, QN => n8017);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           n_1364, QN => n8016);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           n_1365, QN => n8015);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           n_1366, QN => n8014);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           n_1367, QN => n8013);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           n_1368, QN => n8012);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           n_1369, QN => n8011);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           n_1370, QN => n8010);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           n_1371, QN => n8009);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           n_1372, QN => n8008);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           n_1373, QN => n8007);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           n_1374, QN => n8006);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           n_1375, QN => n8005);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           n_1376, QN => n8004);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           n_1377, QN => n8003);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           n_1378, QN => n8002);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           n_1379, QN => n8001);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           n_1380, QN => n8000);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           n_1381, QN => n7999);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           n_1382, QN => n7998);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           n_1383, QN => n7997);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => OUT1_31_port
                           , QN => n_1384);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => OUT1_30_port
                           , QN => n_1385);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => OUT1_29_port
                           , QN => n_1386);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => OUT1_28_port
                           , QN => n_1387);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => OUT1_27_port
                           , QN => n_1388);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => OUT1_26_port
                           , QN => n_1389);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => OUT1_25_port
                           , QN => n_1390);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => OUT1_24_port
                           , QN => n_1391);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => OUT1_23_port
                           , QN => n_1392);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => OUT1_22_port
                           , QN => n_1393);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => OUT1_21_port
                           , QN => n_1394);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => OUT1_20_port
                           , QN => n_1395);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => OUT1_19_port
                           , QN => n_1396);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => OUT1_18_port
                           , QN => n_1397);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => OUT1_17_port
                           , QN => n_1398);
   OUT1_reg_16_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => OUT1_16_port
                           , QN => n_1399);
   OUT1_reg_15_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => OUT1_15_port
                           , QN => n_1400);
   OUT1_reg_14_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => OUT1_14_port
                           , QN => n_1401);
   OUT1_reg_13_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => OUT1_13_port
                           , QN => n_1402);
   OUT1_reg_12_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => OUT1_12_port
                           , QN => n_1403);
   OUT1_reg_11_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => OUT1_11_port
                           , QN => n_1404);
   OUT1_reg_10_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => OUT1_10_port
                           , QN => n_1405);
   OUT1_reg_9_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => OUT1_9_port, 
                           QN => n_1406);
   OUT1_reg_8_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => OUT1_8_port, 
                           QN => n_1407);
   OUT1_reg_7_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1408);
   OUT1_reg_6_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1409);
   OUT1_reg_5_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1410);
   OUT1_reg_4_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1411);
   OUT1_reg_3_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1412);
   OUT1_reg_2_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1413);
   OUT1_reg_1_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1414);
   OUT1_reg_0_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1415);
   OUT2_reg_31_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => OUT2_31_port
                           , QN => n_1416);
   OUT2_reg_30_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => OUT2_30_port
                           , QN => n_1417);
   OUT2_reg_29_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => OUT2_29_port
                           , QN => n_1418);
   OUT2_reg_28_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => OUT2_28_port
                           , QN => n_1419);
   OUT2_reg_27_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => OUT2_27_port
                           , QN => n_1420);
   OUT2_reg_26_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => OUT2_26_port
                           , QN => n_1421);
   OUT2_reg_25_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => OUT2_25_port
                           , QN => n_1422);
   OUT2_reg_24_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => OUT2_24_port
                           , QN => n_1423);
   OUT2_reg_23_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => OUT2_23_port
                           , QN => n_1424);
   OUT2_reg_22_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => OUT2_22_port
                           , QN => n_1425);
   OUT2_reg_21_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => OUT2_21_port
                           , QN => n_1426);
   OUT2_reg_20_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => OUT2_20_port
                           , QN => n_1427);
   OUT2_reg_19_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => OUT2_19_port
                           , QN => n_1428);
   OUT2_reg_18_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => OUT2_18_port
                           , QN => n_1429);
   OUT2_reg_17_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => OUT2_17_port
                           , QN => n_1430);
   OUT2_reg_16_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => OUT2_16_port
                           , QN => n_1431);
   OUT2_reg_15_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => OUT2_15_port
                           , QN => n_1432);
   OUT2_reg_14_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => OUT2_14_port
                           , QN => n_1433);
   OUT2_reg_13_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => OUT2_13_port
                           , QN => n_1434);
   OUT2_reg_12_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => OUT2_12_port
                           , QN => n_1435);
   OUT2_reg_11_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => OUT2_11_port
                           , QN => n_1436);
   OUT2_reg_10_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => OUT2_10_port
                           , QN => n_1437);
   OUT2_reg_9_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1438);
   OUT2_reg_8_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1439);
   OUT2_reg_7_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1440);
   OUT2_reg_6_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1441);
   OUT2_reg_5_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1442);
   OUT2_reg_4_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1443);
   OUT2_reg_3_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1444);
   OUT2_reg_2_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1445);
   OUT2_reg_1_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1446);
   OUT2_reg_0_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1447);
   U3247 : NAND3_X1 port map( A1 => ENABLE, A2 => n9025, A3 => RD2, ZN => n884)
                           ;
   U3248 : NAND3_X1 port map( A1 => ENABLE, A2 => n9025, A3 => RD1, ZN => n2506
                           );
   U3249 : NAND3_X1 port map( A1 => n837, A2 => n836, A3 => n838, ZN => n3149);
   U3250 : NAND3_X1 port map( A1 => n837, A2 => n836, A3 => ADD_WR(0), ZN => 
                           n3151);
   U3251 : NAND3_X1 port map( A1 => n838, A2 => n836, A3 => ADD_WR(1), ZN => 
                           n3153);
   U3252 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n836, A3 => ADD_WR(1), ZN 
                           => n3155);
   U3253 : NAND3_X1 port map( A1 => n838, A2 => n837, A3 => ADD_WR(2), ZN => 
                           n3157);
   U3254 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n837, A3 => ADD_WR(2), ZN 
                           => n3159);
   U3255 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n838, A3 => ADD_WR(2), ZN 
                           => n3161);
   U3256 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n3163);
   U3 : NOR3_X1 port map( A1 => n8957, A2 => ADD_RD2(1), A3 => n848, ZN => 
                           n2473);
   U4 : NOR3_X1 port map( A1 => n8957, A2 => ADD_RD2(0), A3 => n847, ZN => 
                           n2480);
   U5 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n8957, ZN 
                           => n2472);
   U6 : NOR3_X1 port map( A1 => n8909, A2 => ADD_RD1(0), A3 => n842, ZN => 
                           n3095);
   U7 : NOR3_X1 port map( A1 => n847, A2 => n8957, A3 => n848, ZN => n2475);
   U8 : NOR3_X1 port map( A1 => n842, A2 => n8909, A3 => n843, ZN => n3102);
   U9 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n8909, ZN 
                           => n3099);
   U10 : NOR3_X1 port map( A1 => n8909, A2 => ADD_RD1(1), A3 => n843, ZN => 
                           n3096);
   U11 : INV_X1 port map( A => n8454, ZN => n8447);
   U12 : INV_X1 port map( A => n8463, ZN => n8456);
   U13 : INV_X1 port map( A => n8472, ZN => n8465);
   U14 : INV_X1 port map( A => n8481, ZN => n8474);
   U15 : INV_X1 port map( A => n8490, ZN => n8483);
   U16 : INV_X1 port map( A => n8499, ZN => n8492);
   U17 : INV_X1 port map( A => n8508, ZN => n8501);
   U18 : INV_X1 port map( A => n8517, ZN => n8510);
   U19 : INV_X1 port map( A => n8526, ZN => n8519);
   U20 : INV_X1 port map( A => n8535, ZN => n8528);
   U21 : INV_X1 port map( A => n8544, ZN => n8537);
   U22 : INV_X1 port map( A => n8553, ZN => n8546);
   U23 : INV_X1 port map( A => n8562, ZN => n8555);
   U24 : INV_X1 port map( A => n8571, ZN => n8564);
   U25 : INV_X1 port map( A => n8580, ZN => n8573);
   U26 : INV_X1 port map( A => n8589, ZN => n8582);
   U27 : INV_X1 port map( A => n8598, ZN => n8591);
   U28 : INV_X1 port map( A => n8607, ZN => n8600);
   U29 : INV_X1 port map( A => n8616, ZN => n8609);
   U30 : INV_X1 port map( A => n8625, ZN => n8618);
   U31 : INV_X1 port map( A => n8634, ZN => n8627);
   U32 : INV_X1 port map( A => n8643, ZN => n8636);
   U33 : INV_X1 port map( A => n8652, ZN => n8645);
   U34 : INV_X1 port map( A => n8661, ZN => n8654);
   U35 : INV_X1 port map( A => n8670, ZN => n8663);
   U36 : INV_X1 port map( A => n8679, ZN => n8672);
   U37 : INV_X1 port map( A => n8688, ZN => n8681);
   U38 : INV_X1 port map( A => n8697, ZN => n8690);
   U39 : INV_X1 port map( A => n8706, ZN => n8699);
   U40 : INV_X1 port map( A => n8715, ZN => n8708);
   U41 : INV_X1 port map( A => n8817, ZN => n8810);
   U42 : BUF_X1 port map( A => n895, Z => n8931);
   U43 : BUF_X1 port map( A => n895, Z => n8930);
   U44 : BUF_X1 port map( A => n2513, Z => n8892);
   U45 : BUF_X1 port map( A => n2513, Z => n8891);
   U46 : BUF_X1 port map( A => n2517, Z => n8883);
   U47 : BUF_X1 port map( A => n2517, Z => n8882);
   U48 : BUF_X1 port map( A => n895, Z => n8932);
   U49 : BUF_X1 port map( A => n891, Z => n8940);
   U50 : BUF_X1 port map( A => n891, Z => n8939);
   U51 : BUF_X1 port map( A => n2513, Z => n8893);
   U52 : BUF_X1 port map( A => n2517, Z => n8884);
   U53 : BUF_X1 port map( A => n891, Z => n8941);
   U54 : BUF_X1 port map( A => n8446, Z => n8438);
   U55 : BUF_X1 port map( A => n8446, Z => n8439);
   U56 : BUF_X1 port map( A => n8446, Z => n8440);
   U57 : BUF_X1 port map( A => n8446, Z => n8441);
   U58 : BUF_X1 port map( A => n8446, Z => n8442);
   U59 : BUF_X1 port map( A => n8446, Z => n8443);
   U60 : BUF_X1 port map( A => n8443, Z => n8444);
   U61 : BUF_X1 port map( A => n8438, Z => n8445);
   U62 : NAND2_X1 port map( A1 => n2475, A2 => n2471, ZN => n891);
   U63 : BUF_X1 port map( A => n893, Z => n8937);
   U64 : BUF_X1 port map( A => n898, Z => n8925);
   U65 : BUF_X1 port map( A => n858, Z => n9012);
   U66 : BUF_X1 port map( A => n863, Z => n9000);
   U67 : BUF_X1 port map( A => n868, Z => n8988);
   U68 : BUF_X1 port map( A => n893, Z => n8936);
   U69 : BUF_X1 port map( A => n898, Z => n8924);
   U70 : BUF_X1 port map( A => n858, Z => n9011);
   U71 : BUF_X1 port map( A => n863, Z => n8999);
   U72 : BUF_X1 port map( A => n868, Z => n8987);
   U73 : BUF_X1 port map( A => n885, Z => n8955);
   U74 : BUF_X1 port map( A => n880, Z => n8967);
   U75 : BUF_X1 port map( A => n890, Z => n8943);
   U76 : BUF_X1 port map( A => n855, Z => n9018);
   U77 : BUF_X1 port map( A => n885, Z => n8954);
   U78 : BUF_X1 port map( A => n880, Z => n8966);
   U79 : BUF_X1 port map( A => n890, Z => n8942);
   U80 : BUF_X1 port map( A => n855, Z => n9017);
   U81 : BUF_X1 port map( A => n889, Z => n8946);
   U82 : BUF_X1 port map( A => n894, Z => n8934);
   U83 : BUF_X1 port map( A => n899, Z => n8922);
   U84 : BUF_X1 port map( A => n859, Z => n9009);
   U85 : BUF_X1 port map( A => n864, Z => n8997);
   U86 : BUF_X1 port map( A => n869, Z => n8985);
   U87 : BUF_X1 port map( A => n889, Z => n8945);
   U88 : BUF_X1 port map( A => n894, Z => n8933);
   U89 : BUF_X1 port map( A => n899, Z => n8921);
   U90 : BUF_X1 port map( A => n859, Z => n9008);
   U91 : BUF_X1 port map( A => n864, Z => n8996);
   U92 : BUF_X1 port map( A => n869, Z => n8984);
   U93 : BUF_X1 port map( A => n874, Z => n8973);
   U94 : BUF_X1 port map( A => n874, Z => n8972);
   U95 : BUF_X1 port map( A => n2528, Z => n8865);
   U96 : BUF_X1 port map( A => n2526, Z => n8871);
   U97 : BUF_X1 port map( A => n2530, Z => n8859);
   U98 : BUF_X1 port map( A => n2538, Z => n8838);
   U99 : BUF_X1 port map( A => n2543, Z => n8826);
   U100 : BUF_X1 port map( A => n2528, Z => n8864);
   U101 : BUF_X1 port map( A => n2526, Z => n8870);
   U102 : BUF_X1 port map( A => n2530, Z => n8858);
   U103 : BUF_X1 port map( A => n2538, Z => n8837);
   U104 : BUF_X1 port map( A => n2543, Z => n8825);
   U105 : NAND2_X1 port map( A1 => n3102, A2 => n3103, ZN => n2513);
   U106 : BUF_X1 port map( A => n2529, Z => n8862);
   U107 : BUF_X1 port map( A => n2527, Z => n8868);
   U108 : BUF_X1 port map( A => n2531, Z => n8856);
   U109 : BUF_X1 port map( A => n2539, Z => n8835);
   U110 : BUF_X1 port map( A => n2544, Z => n8823);
   U111 : BUF_X1 port map( A => n2529, Z => n8861);
   U112 : BUF_X1 port map( A => n2527, Z => n8867);
   U113 : BUF_X1 port map( A => n2531, Z => n8855);
   U114 : BUF_X1 port map( A => n2539, Z => n8834);
   U115 : BUF_X1 port map( A => n2544, Z => n8822);
   U116 : BUF_X1 port map( A => n875, Z => n8970);
   U117 : BUF_X1 port map( A => n875, Z => n8969);
   U118 : BUF_X1 port map( A => n886, Z => n8952);
   U119 : BUF_X1 port map( A => n881, Z => n8964);
   U120 : BUF_X1 port map( A => n871, Z => n8979);
   U121 : BUF_X1 port map( A => n861, Z => n9003);
   U122 : BUF_X1 port map( A => n866, Z => n8991);
   U123 : BUF_X1 port map( A => n886, Z => n8951);
   U124 : BUF_X1 port map( A => n881, Z => n8963);
   U125 : BUF_X1 port map( A => n871, Z => n8978);
   U126 : BUF_X1 port map( A => n861, Z => n9002);
   U127 : BUF_X1 port map( A => n866, Z => n8990);
   U128 : BUF_X1 port map( A => n2508, Z => n8904);
   U129 : BUF_X1 port map( A => n2503, Z => n8916);
   U130 : BUF_X1 port map( A => n2518, Z => n8880);
   U131 : BUF_X1 port map( A => n2508, Z => n8903);
   U132 : BUF_X1 port map( A => n2503, Z => n8915);
   U133 : BUF_X1 port map( A => n2518, Z => n8879);
   U134 : BUF_X1 port map( A => n2535, Z => n8844);
   U135 : BUF_X1 port map( A => n2540, Z => n8832);
   U136 : BUF_X1 port map( A => n2535, Z => n8843);
   U137 : BUF_X1 port map( A => n2540, Z => n8831);
   U138 : BUF_X1 port map( A => n873, Z => n8976);
   U139 : BUF_X1 port map( A => n873, Z => n8975);
   U140 : BUF_X1 port map( A => n888, Z => n8949);
   U141 : BUF_X1 port map( A => n883, Z => n8961);
   U142 : BUF_X1 port map( A => n888, Z => n8948);
   U143 : BUF_X1 port map( A => n883, Z => n8960);
   U144 : BUF_X1 port map( A => n2510, Z => n8901);
   U145 : BUF_X1 port map( A => n2505, Z => n8913);
   U146 : BUF_X1 port map( A => n2515, Z => n8889);
   U147 : BUF_X1 port map( A => n2520, Z => n8877);
   U148 : BUF_X1 port map( A => n2510, Z => n8900);
   U149 : BUF_X1 port map( A => n2505, Z => n8912);
   U150 : BUF_X1 port map( A => n2515, Z => n8888);
   U151 : BUF_X1 port map( A => n2520, Z => n8876);
   U152 : BUF_X1 port map( A => n2536, Z => n8841);
   U153 : BUF_X1 port map( A => n2541, Z => n8829);
   U154 : BUF_X1 port map( A => n2536, Z => n8840);
   U155 : BUF_X1 port map( A => n2541, Z => n8828);
   U156 : BUF_X1 port map( A => n870, Z => n8982);
   U157 : BUF_X1 port map( A => n860, Z => n9006);
   U158 : BUF_X1 port map( A => n865, Z => n8994);
   U159 : BUF_X1 port map( A => n870, Z => n8981);
   U160 : BUF_X1 port map( A => n860, Z => n9005);
   U161 : BUF_X1 port map( A => n865, Z => n8993);
   U162 : BUF_X1 port map( A => n2507, Z => n8907);
   U163 : BUF_X1 port map( A => n2502, Z => n8919);
   U164 : BUF_X1 port map( A => n2512, Z => n8895);
   U165 : BUF_X1 port map( A => n2507, Z => n8906);
   U166 : BUF_X1 port map( A => n2502, Z => n8918);
   U167 : BUF_X1 port map( A => n2512, Z => n8894);
   U168 : BUF_X1 port map( A => n893, Z => n8938);
   U169 : BUF_X1 port map( A => n898, Z => n8926);
   U170 : BUF_X1 port map( A => n858, Z => n9013);
   U171 : BUF_X1 port map( A => n863, Z => n9001);
   U172 : BUF_X1 port map( A => n868, Z => n8989);
   U173 : BUF_X1 port map( A => n885, Z => n8956);
   U174 : BUF_X1 port map( A => n880, Z => n8968);
   U175 : BUF_X1 port map( A => n890, Z => n8944);
   U176 : BUF_X1 port map( A => n855, Z => n9019);
   U177 : BUF_X1 port map( A => n899, Z => n8923);
   U178 : BUF_X1 port map( A => n889, Z => n8947);
   U179 : BUF_X1 port map( A => n894, Z => n8935);
   U180 : BUF_X1 port map( A => n859, Z => n9010);
   U181 : BUF_X1 port map( A => n864, Z => n8998);
   U182 : BUF_X1 port map( A => n869, Z => n8986);
   U183 : BUF_X1 port map( A => n2534, Z => n8847);
   U184 : BUF_X1 port map( A => n2534, Z => n8846);
   U185 : BUF_X1 port map( A => n874, Z => n8974);
   U186 : BUF_X1 port map( A => n2528, Z => n8866);
   U187 : BUF_X1 port map( A => n2526, Z => n8872);
   U188 : BUF_X1 port map( A => n2530, Z => n8860);
   U189 : BUF_X1 port map( A => n2538, Z => n8839);
   U190 : BUF_X1 port map( A => n2543, Z => n8827);
   U191 : BUF_X1 port map( A => n2532, Z => n8853);
   U192 : BUF_X1 port map( A => n2532, Z => n8852);
   U193 : BUF_X1 port map( A => n2533, Z => n8850);
   U194 : BUF_X1 port map( A => n2533, Z => n8849);
   U195 : BUF_X1 port map( A => n896, Z => n8928);
   U196 : BUF_X1 port map( A => n856, Z => n9015);
   U197 : BUF_X1 port map( A => n896, Z => n8927);
   U198 : BUF_X1 port map( A => n856, Z => n9014);
   U199 : BUF_X1 port map( A => n2529, Z => n8863);
   U200 : BUF_X1 port map( A => n2527, Z => n8869);
   U201 : BUF_X1 port map( A => n2531, Z => n8857);
   U202 : BUF_X1 port map( A => n2539, Z => n8836);
   U203 : BUF_X1 port map( A => n2544, Z => n8824);
   U204 : BUF_X1 port map( A => n2511, Z => n8897);
   U205 : BUF_X1 port map( A => n2516, Z => n8885);
   U206 : BUF_X1 port map( A => n2521, Z => n8873);
   U207 : BUF_X1 port map( A => n2511, Z => n8898);
   U208 : BUF_X1 port map( A => n2516, Z => n8886);
   U209 : BUF_X1 port map( A => n2521, Z => n8874);
   U210 : BUF_X1 port map( A => n875, Z => n8971);
   U211 : BUF_X1 port map( A => n886, Z => n8953);
   U212 : BUF_X1 port map( A => n881, Z => n8965);
   U213 : BUF_X1 port map( A => n871, Z => n8980);
   U214 : BUF_X1 port map( A => n861, Z => n9004);
   U215 : BUF_X1 port map( A => n866, Z => n8992);
   U216 : BUF_X1 port map( A => n2508, Z => n8905);
   U217 : BUF_X1 port map( A => n2503, Z => n8917);
   U218 : BUF_X1 port map( A => n2518, Z => n8881);
   U219 : BUF_X1 port map( A => n2535, Z => n8845);
   U220 : BUF_X1 port map( A => n2540, Z => n8833);
   U221 : BUF_X1 port map( A => n873, Z => n8977);
   U222 : BUF_X1 port map( A => n888, Z => n8950);
   U223 : BUF_X1 port map( A => n883, Z => n8962);
   U224 : BUF_X1 port map( A => n2510, Z => n8902);
   U225 : BUF_X1 port map( A => n2505, Z => n8914);
   U226 : BUF_X1 port map( A => n2515, Z => n8890);
   U227 : BUF_X1 port map( A => n2520, Z => n8878);
   U228 : BUF_X1 port map( A => n2541, Z => n8830);
   U229 : BUF_X1 port map( A => n2536, Z => n8842);
   U230 : BUF_X1 port map( A => n870, Z => n8983);
   U231 : BUF_X1 port map( A => n860, Z => n9007);
   U232 : BUF_X1 port map( A => n865, Z => n8995);
   U233 : BUF_X1 port map( A => n2507, Z => n8908);
   U234 : BUF_X1 port map( A => n2502, Z => n8920);
   U235 : BUF_X1 port map( A => n2512, Z => n8896);
   U236 : BUF_X1 port map( A => n2534, Z => n8848);
   U237 : BUF_X1 port map( A => n2532, Z => n8854);
   U238 : BUF_X1 port map( A => n2533, Z => n8851);
   U239 : BUF_X1 port map( A => n896, Z => n8929);
   U240 : BUF_X1 port map( A => n856, Z => n9016);
   U241 : BUF_X1 port map( A => n2511, Z => n8899);
   U242 : BUF_X1 port map( A => n2516, Z => n8887);
   U243 : BUF_X1 port map( A => n2521, Z => n8875);
   U244 : NAND2_X1 port map( A1 => n2489, A2 => n2475, ZN => n895);
   U245 : NAND2_X1 port map( A1 => n3094, A2 => n3102, ZN => n2517);
   U246 : BUF_X1 port map( A => n8455, Z => n8448);
   U247 : BUF_X1 port map( A => n8455, Z => n8449);
   U248 : BUF_X1 port map( A => n8455, Z => n8450);
   U249 : BUF_X1 port map( A => n8455, Z => n8451);
   U250 : BUF_X1 port map( A => n8455, Z => n8452);
   U251 : BUF_X1 port map( A => n8455, Z => n8453);
   U252 : BUF_X1 port map( A => n8464, Z => n8457);
   U253 : BUF_X1 port map( A => n8464, Z => n8458);
   U254 : BUF_X1 port map( A => n8464, Z => n8459);
   U255 : BUF_X1 port map( A => n8464, Z => n8460);
   U256 : BUF_X1 port map( A => n8464, Z => n8461);
   U257 : BUF_X1 port map( A => n8464, Z => n8462);
   U258 : BUF_X1 port map( A => n8473, Z => n8466);
   U259 : BUF_X1 port map( A => n8473, Z => n8467);
   U260 : BUF_X1 port map( A => n8473, Z => n8468);
   U261 : BUF_X1 port map( A => n8473, Z => n8469);
   U262 : BUF_X1 port map( A => n8473, Z => n8470);
   U263 : BUF_X1 port map( A => n8473, Z => n8471);
   U264 : BUF_X1 port map( A => n8482, Z => n8475);
   U265 : BUF_X1 port map( A => n8482, Z => n8476);
   U266 : BUF_X1 port map( A => n8482, Z => n8477);
   U267 : BUF_X1 port map( A => n8482, Z => n8478);
   U268 : BUF_X1 port map( A => n8482, Z => n8479);
   U269 : BUF_X1 port map( A => n8482, Z => n8480);
   U270 : BUF_X1 port map( A => n8491, Z => n8484);
   U271 : BUF_X1 port map( A => n8491, Z => n8485);
   U272 : BUF_X1 port map( A => n8491, Z => n8486);
   U273 : BUF_X1 port map( A => n8491, Z => n8487);
   U274 : BUF_X1 port map( A => n8491, Z => n8488);
   U275 : BUF_X1 port map( A => n8491, Z => n8489);
   U276 : BUF_X1 port map( A => n8500, Z => n8493);
   U277 : BUF_X1 port map( A => n8500, Z => n8494);
   U278 : BUF_X1 port map( A => n8500, Z => n8495);
   U279 : BUF_X1 port map( A => n8500, Z => n8496);
   U280 : BUF_X1 port map( A => n8500, Z => n8497);
   U281 : BUF_X1 port map( A => n8500, Z => n8498);
   U282 : BUF_X1 port map( A => n8509, Z => n8502);
   U283 : BUF_X1 port map( A => n8509, Z => n8503);
   U284 : BUF_X1 port map( A => n8509, Z => n8504);
   U285 : BUF_X1 port map( A => n8509, Z => n8505);
   U286 : BUF_X1 port map( A => n8509, Z => n8506);
   U287 : BUF_X1 port map( A => n8509, Z => n8507);
   U288 : BUF_X1 port map( A => n8518, Z => n8511);
   U289 : BUF_X1 port map( A => n8518, Z => n8512);
   U290 : BUF_X1 port map( A => n8518, Z => n8513);
   U291 : BUF_X1 port map( A => n8518, Z => n8514);
   U292 : BUF_X1 port map( A => n8518, Z => n8515);
   U293 : BUF_X1 port map( A => n8518, Z => n8516);
   U294 : BUF_X1 port map( A => n8527, Z => n8520);
   U295 : BUF_X1 port map( A => n8527, Z => n8521);
   U296 : BUF_X1 port map( A => n8527, Z => n8522);
   U297 : BUF_X1 port map( A => n8527, Z => n8523);
   U298 : BUF_X1 port map( A => n8527, Z => n8524);
   U299 : BUF_X1 port map( A => n8527, Z => n8525);
   U300 : BUF_X1 port map( A => n8536, Z => n8529);
   U301 : BUF_X1 port map( A => n8536, Z => n8530);
   U302 : BUF_X1 port map( A => n8536, Z => n8531);
   U303 : BUF_X1 port map( A => n8536, Z => n8532);
   U304 : BUF_X1 port map( A => n8536, Z => n8533);
   U305 : BUF_X1 port map( A => n8536, Z => n8534);
   U306 : BUF_X1 port map( A => n8545, Z => n8538);
   U307 : BUF_X1 port map( A => n8545, Z => n8539);
   U308 : BUF_X1 port map( A => n8545, Z => n8540);
   U309 : BUF_X1 port map( A => n8545, Z => n8541);
   U310 : BUF_X1 port map( A => n8545, Z => n8542);
   U311 : BUF_X1 port map( A => n8545, Z => n8543);
   U312 : BUF_X1 port map( A => n8554, Z => n8547);
   U313 : BUF_X1 port map( A => n8554, Z => n8548);
   U314 : BUF_X1 port map( A => n8554, Z => n8549);
   U315 : BUF_X1 port map( A => n8554, Z => n8550);
   U316 : BUF_X1 port map( A => n8554, Z => n8551);
   U317 : BUF_X1 port map( A => n8554, Z => n8552);
   U318 : BUF_X1 port map( A => n8563, Z => n8556);
   U319 : BUF_X1 port map( A => n8563, Z => n8557);
   U320 : BUF_X1 port map( A => n8563, Z => n8558);
   U321 : BUF_X1 port map( A => n8563, Z => n8559);
   U322 : BUF_X1 port map( A => n8563, Z => n8560);
   U323 : BUF_X1 port map( A => n8563, Z => n8561);
   U324 : BUF_X1 port map( A => n8572, Z => n8565);
   U325 : BUF_X1 port map( A => n8572, Z => n8566);
   U326 : BUF_X1 port map( A => n8572, Z => n8567);
   U327 : BUF_X1 port map( A => n8572, Z => n8568);
   U328 : BUF_X1 port map( A => n8572, Z => n8569);
   U329 : BUF_X1 port map( A => n8572, Z => n8570);
   U330 : BUF_X1 port map( A => n8581, Z => n8574);
   U331 : BUF_X1 port map( A => n8581, Z => n8575);
   U332 : BUF_X1 port map( A => n8581, Z => n8576);
   U333 : BUF_X1 port map( A => n8581, Z => n8577);
   U334 : BUF_X1 port map( A => n8581, Z => n8578);
   U335 : BUF_X1 port map( A => n8581, Z => n8579);
   U336 : BUF_X1 port map( A => n8590, Z => n8583);
   U337 : BUF_X1 port map( A => n8590, Z => n8584);
   U338 : BUF_X1 port map( A => n8590, Z => n8585);
   U339 : BUF_X1 port map( A => n8590, Z => n8586);
   U340 : BUF_X1 port map( A => n8590, Z => n8587);
   U341 : BUF_X1 port map( A => n8590, Z => n8588);
   U342 : BUF_X1 port map( A => n8599, Z => n8592);
   U343 : BUF_X1 port map( A => n8599, Z => n8593);
   U344 : BUF_X1 port map( A => n8599, Z => n8594);
   U345 : BUF_X1 port map( A => n8599, Z => n8595);
   U346 : BUF_X1 port map( A => n8599, Z => n8596);
   U347 : BUF_X1 port map( A => n8599, Z => n8597);
   U348 : BUF_X1 port map( A => n8608, Z => n8601);
   U349 : BUF_X1 port map( A => n8608, Z => n8602);
   U350 : BUF_X1 port map( A => n8608, Z => n8603);
   U351 : BUF_X1 port map( A => n8608, Z => n8604);
   U352 : BUF_X1 port map( A => n8608, Z => n8605);
   U353 : BUF_X1 port map( A => n8608, Z => n8606);
   U354 : BUF_X1 port map( A => n8617, Z => n8610);
   U355 : BUF_X1 port map( A => n8617, Z => n8611);
   U356 : BUF_X1 port map( A => n8617, Z => n8612);
   U357 : BUF_X1 port map( A => n8617, Z => n8613);
   U358 : BUF_X1 port map( A => n8617, Z => n8614);
   U359 : BUF_X1 port map( A => n8617, Z => n8615);
   U360 : BUF_X1 port map( A => n8626, Z => n8619);
   U361 : BUF_X1 port map( A => n8626, Z => n8620);
   U362 : BUF_X1 port map( A => n8626, Z => n8621);
   U363 : BUF_X1 port map( A => n8626, Z => n8622);
   U364 : BUF_X1 port map( A => n8626, Z => n8623);
   U365 : BUF_X1 port map( A => n8626, Z => n8624);
   U366 : BUF_X1 port map( A => n8635, Z => n8628);
   U367 : BUF_X1 port map( A => n8635, Z => n8629);
   U368 : BUF_X1 port map( A => n8635, Z => n8630);
   U369 : BUF_X1 port map( A => n8635, Z => n8631);
   U370 : BUF_X1 port map( A => n8635, Z => n8632);
   U371 : BUF_X1 port map( A => n8635, Z => n8633);
   U372 : BUF_X1 port map( A => n8644, Z => n8637);
   U373 : BUF_X1 port map( A => n8644, Z => n8638);
   U374 : BUF_X1 port map( A => n8644, Z => n8639);
   U375 : BUF_X1 port map( A => n8644, Z => n8640);
   U376 : BUF_X1 port map( A => n8644, Z => n8641);
   U377 : BUF_X1 port map( A => n8644, Z => n8642);
   U378 : BUF_X1 port map( A => n8653, Z => n8646);
   U379 : BUF_X1 port map( A => n8653, Z => n8647);
   U380 : BUF_X1 port map( A => n8653, Z => n8648);
   U381 : BUF_X1 port map( A => n8653, Z => n8649);
   U382 : BUF_X1 port map( A => n8653, Z => n8650);
   U383 : BUF_X1 port map( A => n8653, Z => n8651);
   U384 : BUF_X1 port map( A => n8662, Z => n8655);
   U385 : BUF_X1 port map( A => n8662, Z => n8656);
   U386 : BUF_X1 port map( A => n8662, Z => n8657);
   U387 : BUF_X1 port map( A => n8662, Z => n8658);
   U388 : BUF_X1 port map( A => n8662, Z => n8659);
   U389 : BUF_X1 port map( A => n8662, Z => n8660);
   U390 : BUF_X1 port map( A => n8671, Z => n8664);
   U391 : BUF_X1 port map( A => n8671, Z => n8665);
   U392 : BUF_X1 port map( A => n8671, Z => n8666);
   U393 : BUF_X1 port map( A => n8671, Z => n8667);
   U394 : BUF_X1 port map( A => n8671, Z => n8668);
   U395 : BUF_X1 port map( A => n8671, Z => n8669);
   U396 : BUF_X1 port map( A => n8680, Z => n8673);
   U397 : BUF_X1 port map( A => n8680, Z => n8674);
   U398 : BUF_X1 port map( A => n8680, Z => n8675);
   U399 : BUF_X1 port map( A => n8680, Z => n8676);
   U400 : BUF_X1 port map( A => n8680, Z => n8677);
   U401 : BUF_X1 port map( A => n8680, Z => n8678);
   U402 : BUF_X1 port map( A => n8689, Z => n8682);
   U403 : BUF_X1 port map( A => n8689, Z => n8683);
   U404 : BUF_X1 port map( A => n8689, Z => n8684);
   U405 : BUF_X1 port map( A => n8689, Z => n8685);
   U406 : BUF_X1 port map( A => n8689, Z => n8686);
   U407 : BUF_X1 port map( A => n8689, Z => n8687);
   U408 : BUF_X1 port map( A => n8698, Z => n8691);
   U409 : BUF_X1 port map( A => n8698, Z => n8692);
   U410 : BUF_X1 port map( A => n8698, Z => n8693);
   U411 : BUF_X1 port map( A => n8698, Z => n8694);
   U412 : BUF_X1 port map( A => n8698, Z => n8695);
   U413 : BUF_X1 port map( A => n8698, Z => n8696);
   U414 : BUF_X1 port map( A => n8707, Z => n8700);
   U415 : BUF_X1 port map( A => n8707, Z => n8701);
   U416 : BUF_X1 port map( A => n8707, Z => n8702);
   U417 : BUF_X1 port map( A => n8707, Z => n8703);
   U418 : BUF_X1 port map( A => n8707, Z => n8704);
   U419 : BUF_X1 port map( A => n8707, Z => n8705);
   U420 : BUF_X1 port map( A => n8716, Z => n8709);
   U421 : BUF_X1 port map( A => n8716, Z => n8710);
   U422 : BUF_X1 port map( A => n8716, Z => n8711);
   U423 : BUF_X1 port map( A => n8716, Z => n8712);
   U424 : BUF_X1 port map( A => n8716, Z => n8713);
   U425 : BUF_X1 port map( A => n8716, Z => n8714);
   U426 : BUF_X1 port map( A => n8818, Z => n8811);
   U427 : BUF_X1 port map( A => n8818, Z => n8812);
   U428 : BUF_X1 port map( A => n8818, Z => n8813);
   U429 : BUF_X1 port map( A => n8818, Z => n8814);
   U430 : BUF_X1 port map( A => n8818, Z => n8815);
   U431 : BUF_X1 port map( A => n8818, Z => n8816);
   U432 : BUF_X1 port map( A => n8455, Z => n8454);
   U433 : BUF_X1 port map( A => n8464, Z => n8463);
   U434 : BUF_X1 port map( A => n8473, Z => n8472);
   U435 : BUF_X1 port map( A => n8482, Z => n8481);
   U436 : BUF_X1 port map( A => n8491, Z => n8490);
   U437 : BUF_X1 port map( A => n8500, Z => n8499);
   U438 : BUF_X1 port map( A => n8509, Z => n8508);
   U439 : BUF_X1 port map( A => n8518, Z => n8517);
   U440 : BUF_X1 port map( A => n8527, Z => n8526);
   U441 : BUF_X1 port map( A => n8536, Z => n8535);
   U442 : BUF_X1 port map( A => n8545, Z => n8544);
   U443 : BUF_X1 port map( A => n8554, Z => n8553);
   U444 : BUF_X1 port map( A => n8563, Z => n8562);
   U445 : BUF_X1 port map( A => n8572, Z => n8571);
   U446 : BUF_X1 port map( A => n8581, Z => n8580);
   U447 : BUF_X1 port map( A => n8590, Z => n8589);
   U448 : BUF_X1 port map( A => n8599, Z => n8598);
   U449 : BUF_X1 port map( A => n8608, Z => n8607);
   U450 : BUF_X1 port map( A => n8617, Z => n8616);
   U451 : BUF_X1 port map( A => n8626, Z => n8625);
   U452 : BUF_X1 port map( A => n8635, Z => n8634);
   U453 : BUF_X1 port map( A => n8644, Z => n8643);
   U454 : BUF_X1 port map( A => n8653, Z => n8652);
   U455 : BUF_X1 port map( A => n8662, Z => n8661);
   U456 : BUF_X1 port map( A => n8671, Z => n8670);
   U457 : BUF_X1 port map( A => n8680, Z => n8679);
   U458 : BUF_X1 port map( A => n8689, Z => n8688);
   U459 : BUF_X1 port map( A => n8698, Z => n8697);
   U460 : BUF_X1 port map( A => n8707, Z => n8706);
   U461 : BUF_X1 port map( A => n8716, Z => n8715);
   U462 : BUF_X1 port map( A => n8818, Z => n8817);
   U463 : INV_X1 port map( A => n8437, ZN => n8446);
   U464 : OAI222_X1 port map( A1 => n8181, A2 => n8854, B1 => n7729, B2 => 
                           n8851, C1 => n7889, C2 => n8848, ZN => n2522);
   U465 : OAI222_X1 port map( A1 => n8182, A2 => n8854, B1 => n7730, B2 => 
                           n8851, C1 => n7890, C2 => n8848, ZN => n2557);
   U466 : OAI222_X1 port map( A1 => n8183, A2 => n8854, B1 => n7731, B2 => 
                           n8851, C1 => n7891, C2 => n8848, ZN => n2575);
   U467 : OAI222_X1 port map( A1 => n8184, A2 => n8854, B1 => n7732, B2 => 
                           n8851, C1 => n7892, C2 => n8848, ZN => n2593);
   U468 : OAI222_X1 port map( A1 => n8185, A2 => n8854, B1 => n7733, B2 => 
                           n8851, C1 => n7893, C2 => n8848, ZN => n2611);
   U469 : OAI222_X1 port map( A1 => n8186, A2 => n8854, B1 => n7734, B2 => 
                           n8851, C1 => n7894, C2 => n8848, ZN => n2629);
   U470 : OAI222_X1 port map( A1 => n8187, A2 => n8854, B1 => n7735, B2 => 
                           n8851, C1 => n7895, C2 => n8848, ZN => n2647);
   U471 : OAI222_X1 port map( A1 => n8188, A2 => n8854, B1 => n7736, B2 => 
                           n8851, C1 => n7896, C2 => n8848, ZN => n2665);
   U472 : OAI222_X1 port map( A1 => n8189, A2 => n8853, B1 => n7737, B2 => 
                           n8850, C1 => n7897, C2 => n8847, ZN => n2683);
   U473 : OAI222_X1 port map( A1 => n8190, A2 => n8853, B1 => n7738, B2 => 
                           n8850, C1 => n7898, C2 => n8847, ZN => n2701);
   U474 : OAI222_X1 port map( A1 => n8191, A2 => n8853, B1 => n7739, B2 => 
                           n8850, C1 => n7899, C2 => n8847, ZN => n2719);
   U475 : OAI222_X1 port map( A1 => n8192, A2 => n8853, B1 => n7740, B2 => 
                           n8850, C1 => n7900, C2 => n8847, ZN => n2737);
   U476 : OAI222_X1 port map( A1 => n8193, A2 => n8853, B1 => n7645, B2 => 
                           n8850, C1 => n7769, C2 => n8847, ZN => n2755);
   U477 : OAI222_X1 port map( A1 => n8194, A2 => n8853, B1 => n7646, B2 => 
                           n8850, C1 => n7770, C2 => n8847, ZN => n2773);
   U478 : OAI222_X1 port map( A1 => n8195, A2 => n8853, B1 => n7647, B2 => 
                           n8850, C1 => n7771, C2 => n8847, ZN => n2791);
   U479 : OAI222_X1 port map( A1 => n8196, A2 => n8853, B1 => n7648, B2 => 
                           n8850, C1 => n7772, C2 => n8847, ZN => n2809);
   U480 : OAI222_X1 port map( A1 => n8197, A2 => n8853, B1 => n7649, B2 => 
                           n8850, C1 => n7773, C2 => n8847, ZN => n2827);
   U481 : OAI222_X1 port map( A1 => n8198, A2 => n8853, B1 => n7650, B2 => 
                           n8850, C1 => n7774, C2 => n8847, ZN => n2845);
   U482 : OAI222_X1 port map( A1 => n8199, A2 => n8853, B1 => n7651, B2 => 
                           n8850, C1 => n7775, C2 => n8847, ZN => n2863);
   U483 : OAI222_X1 port map( A1 => n8200, A2 => n8853, B1 => n7652, B2 => 
                           n8850, C1 => n7776, C2 => n8847, ZN => n2881);
   U484 : OAI222_X1 port map( A1 => n8201, A2 => n8852, B1 => n7653, B2 => 
                           n8849, C1 => n7777, C2 => n8846, ZN => n2899);
   U485 : OAI222_X1 port map( A1 => n8202, A2 => n8852, B1 => n7654, B2 => 
                           n8849, C1 => n7778, C2 => n8846, ZN => n2917);
   U486 : OAI222_X1 port map( A1 => n8203, A2 => n8852, B1 => n7655, B2 => 
                           n8849, C1 => n7779, C2 => n8846, ZN => n2935);
   U487 : OAI222_X1 port map( A1 => n8204, A2 => n8852, B1 => n7656, B2 => 
                           n8849, C1 => n7780, C2 => n8846, ZN => n2953);
   U488 : OAI222_X1 port map( A1 => n7909, A2 => n8852, B1 => n7637, B2 => 
                           n8849, C1 => n7761, C2 => n8846, ZN => n2971);
   U489 : OAI222_X1 port map( A1 => n7910, A2 => n8852, B1 => n7638, B2 => 
                           n8849, C1 => n7762, C2 => n8846, ZN => n2989);
   U490 : OAI222_X1 port map( A1 => n7911, A2 => n8852, B1 => n7639, B2 => 
                           n8849, C1 => n7763, C2 => n8846, ZN => n3007);
   U491 : OAI222_X1 port map( A1 => n7912, A2 => n8852, B1 => n7640, B2 => 
                           n8849, C1 => n7764, C2 => n8846, ZN => n3025);
   U492 : OAI222_X1 port map( A1 => n7913, A2 => n8852, B1 => n7641, B2 => 
                           n8849, C1 => n7765, C2 => n8846, ZN => n3043);
   U493 : OAI222_X1 port map( A1 => n7914, A2 => n8852, B1 => n7642, B2 => 
                           n8849, C1 => n7766, C2 => n8846, ZN => n3061);
   U494 : OAI222_X1 port map( A1 => n7915, A2 => n8852, B1 => n7643, B2 => 
                           n8849, C1 => n7767, C2 => n8846, ZN => n3079);
   U495 : OAI222_X1 port map( A1 => n7916, A2 => n8852, B1 => n7644, B2 => 
                           n8849, C1 => n7768, C2 => n8846, ZN => n3108);
   U496 : OAI22_X1 port map( A1 => n7841, A2 => n8866, B1 => n8109, B2 => n8863
                           , ZN => n2524);
   U497 : OAI22_X1 port map( A1 => n7842, A2 => n8866, B1 => n8110, B2 => n8863
                           , ZN => n2559);
   U498 : OAI22_X1 port map( A1 => n7843, A2 => n8866, B1 => n8111, B2 => n8863
                           , ZN => n2577);
   U499 : OAI22_X1 port map( A1 => n7844, A2 => n8866, B1 => n8112, B2 => n8863
                           , ZN => n2595);
   U500 : OAI22_X1 port map( A1 => n7845, A2 => n8866, B1 => n8113, B2 => n8863
                           , ZN => n2613);
   U501 : OAI22_X1 port map( A1 => n7846, A2 => n8866, B1 => n8114, B2 => n8863
                           , ZN => n2631);
   U502 : OAI22_X1 port map( A1 => n7847, A2 => n8866, B1 => n8115, B2 => n8863
                           , ZN => n2649);
   U503 : OAI22_X1 port map( A1 => n7848, A2 => n8866, B1 => n8116, B2 => n8863
                           , ZN => n2667);
   U504 : OAI22_X1 port map( A1 => n7829, A2 => n8839, B1 => n8085, B2 => n8836
                           , ZN => n2537);
   U505 : OAI22_X1 port map( A1 => n7830, A2 => n8839, B1 => n8086, B2 => n8836
                           , ZN => n2561);
   U506 : OAI22_X1 port map( A1 => n7831, A2 => n8839, B1 => n8087, B2 => n8836
                           , ZN => n2579);
   U507 : OAI22_X1 port map( A1 => n7832, A2 => n8839, B1 => n8088, B2 => n8836
                           , ZN => n2597);
   U508 : OAI22_X1 port map( A1 => n7833, A2 => n8839, B1 => n8089, B2 => n8836
                           , ZN => n2615);
   U509 : OAI22_X1 port map( A1 => n7834, A2 => n8839, B1 => n8090, B2 => n8836
                           , ZN => n2633);
   U510 : OAI22_X1 port map( A1 => n7835, A2 => n8839, B1 => n8091, B2 => n8836
                           , ZN => n2651);
   U511 : OAI22_X1 port map( A1 => n7836, A2 => n8839, B1 => n8092, B2 => n8836
                           , ZN => n2669);
   U512 : OAI22_X1 port map( A1 => n7849, A2 => n8865, B1 => n8117, B2 => n8862
                           , ZN => n2685);
   U513 : OAI22_X1 port map( A1 => n7850, A2 => n8865, B1 => n8118, B2 => n8862
                           , ZN => n2703);
   U514 : OAI22_X1 port map( A1 => n7851, A2 => n8865, B1 => n8119, B2 => n8862
                           , ZN => n2721);
   U515 : OAI22_X1 port map( A1 => n7852, A2 => n8865, B1 => n8120, B2 => n8862
                           , ZN => n2739);
   U516 : OAI22_X1 port map( A1 => n7717, A2 => n8865, B1 => n8121, B2 => n8862
                           , ZN => n2757);
   U517 : OAI22_X1 port map( A1 => n7718, A2 => n8865, B1 => n8122, B2 => n8862
                           , ZN => n2775);
   U518 : OAI22_X1 port map( A1 => n7719, A2 => n8865, B1 => n8123, B2 => n8862
                           , ZN => n2793);
   U519 : OAI22_X1 port map( A1 => n7720, A2 => n8865, B1 => n8124, B2 => n8862
                           , ZN => n2811);
   U520 : OAI22_X1 port map( A1 => n7721, A2 => n8865, B1 => n8125, B2 => n8862
                           , ZN => n2829);
   U521 : OAI22_X1 port map( A1 => n7722, A2 => n8865, B1 => n8126, B2 => n8862
                           , ZN => n2847);
   U522 : OAI22_X1 port map( A1 => n7723, A2 => n8865, B1 => n8127, B2 => n8862
                           , ZN => n2865);
   U523 : OAI22_X1 port map( A1 => n7724, A2 => n8865, B1 => n8128, B2 => n8862
                           , ZN => n2883);
   U524 : OAI22_X1 port map( A1 => n7725, A2 => n8864, B1 => n8129, B2 => n8861
                           , ZN => n2901);
   U525 : OAI22_X1 port map( A1 => n7726, A2 => n8864, B1 => n8130, B2 => n8861
                           , ZN => n2919);
   U526 : OAI22_X1 port map( A1 => n7727, A2 => n8864, B1 => n8131, B2 => n8861
                           , ZN => n2937);
   U527 : OAI22_X1 port map( A1 => n7728, A2 => n8864, B1 => n8132, B2 => n8861
                           , ZN => n2955);
   U528 : OAI22_X1 port map( A1 => n7697, A2 => n8864, B1 => n7861, B2 => n8861
                           , ZN => n2973);
   U529 : OAI22_X1 port map( A1 => n7698, A2 => n8864, B1 => n7862, B2 => n8861
                           , ZN => n2991);
   U530 : OAI22_X1 port map( A1 => n7699, A2 => n8864, B1 => n7863, B2 => n8861
                           , ZN => n3009);
   U531 : OAI22_X1 port map( A1 => n7700, A2 => n8864, B1 => n7864, B2 => n8861
                           , ZN => n3027);
   U532 : OAI22_X1 port map( A1 => n7701, A2 => n8864, B1 => n7865, B2 => n8861
                           , ZN => n3045);
   U533 : OAI22_X1 port map( A1 => n7702, A2 => n8864, B1 => n7866, B2 => n8861
                           , ZN => n3063);
   U534 : OAI22_X1 port map( A1 => n7703, A2 => n8864, B1 => n7867, B2 => n8861
                           , ZN => n3081);
   U535 : OAI22_X1 port map( A1 => n7704, A2 => n8864, B1 => n7868, B2 => n8861
                           , ZN => n3110);
   U536 : OAI22_X1 port map( A1 => n7837, A2 => n8838, B1 => n8093, B2 => n8835
                           , ZN => n2687);
   U537 : OAI22_X1 port map( A1 => n7838, A2 => n8838, B1 => n8094, B2 => n8835
                           , ZN => n2705);
   U538 : OAI22_X1 port map( A1 => n7839, A2 => n8838, B1 => n8095, B2 => n8835
                           , ZN => n2723);
   U539 : OAI22_X1 port map( A1 => n7840, A2 => n8838, B1 => n8096, B2 => n8835
                           , ZN => n2741);
   U540 : OAI22_X1 port map( A1 => n7705, A2 => n8838, B1 => n8097, B2 => n8835
                           , ZN => n2759);
   U541 : OAI22_X1 port map( A1 => n7706, A2 => n8838, B1 => n8098, B2 => n8835
                           , ZN => n2777);
   U542 : OAI22_X1 port map( A1 => n7707, A2 => n8838, B1 => n8099, B2 => n8835
                           , ZN => n2795);
   U543 : OAI22_X1 port map( A1 => n7708, A2 => n8838, B1 => n8100, B2 => n8835
                           , ZN => n2813);
   U544 : OAI22_X1 port map( A1 => n7709, A2 => n8838, B1 => n8101, B2 => n8835
                           , ZN => n2831);
   U545 : OAI22_X1 port map( A1 => n7710, A2 => n8838, B1 => n8102, B2 => n8835
                           , ZN => n2849);
   U546 : OAI22_X1 port map( A1 => n7711, A2 => n8838, B1 => n8103, B2 => n8835
                           , ZN => n2867);
   U547 : OAI22_X1 port map( A1 => n7712, A2 => n8838, B1 => n8104, B2 => n8835
                           , ZN => n2885);
   U548 : OAI22_X1 port map( A1 => n7713, A2 => n8837, B1 => n8105, B2 => n8834
                           , ZN => n2903);
   U549 : OAI22_X1 port map( A1 => n7714, A2 => n8837, B1 => n8106, B2 => n8834
                           , ZN => n2921);
   U550 : OAI22_X1 port map( A1 => n7715, A2 => n8837, B1 => n8107, B2 => n8834
                           , ZN => n2939);
   U551 : OAI22_X1 port map( A1 => n7716, A2 => n8837, B1 => n8108, B2 => n8834
                           , ZN => n2957);
   U552 : OAI22_X1 port map( A1 => n7689, A2 => n8837, B1 => n7853, B2 => n8834
                           , ZN => n2975);
   U553 : OAI22_X1 port map( A1 => n7690, A2 => n8837, B1 => n7854, B2 => n8834
                           , ZN => n2993);
   U554 : OAI22_X1 port map( A1 => n7691, A2 => n8837, B1 => n7855, B2 => n8834
                           , ZN => n3011);
   U555 : OAI22_X1 port map( A1 => n7692, A2 => n8837, B1 => n7856, B2 => n8834
                           , ZN => n3029);
   U556 : OAI22_X1 port map( A1 => n7693, A2 => n8837, B1 => n7857, B2 => n8834
                           , ZN => n3047);
   U557 : OAI22_X1 port map( A1 => n7694, A2 => n8837, B1 => n7858, B2 => n8834
                           , ZN => n3065);
   U558 : OAI22_X1 port map( A1 => n7695, A2 => n8837, B1 => n7859, B2 => n8834
                           , ZN => n3083);
   U559 : OAI22_X1 port map( A1 => n7696, A2 => n8837, B1 => n7860, B2 => n8834
                           , ZN => n3113);
   U560 : OAI22_X1 port map( A1 => n8479, A2 => n8791, B1 => n7821, B2 => n3186
                           , ZN => n1424);
   U561 : OAI22_X1 port map( A1 => n8480, A2 => n8794, B1 => n7822, B2 => n3186
                           , ZN => n1425);
   U562 : OAI22_X1 port map( A1 => n8480, A2 => n8797, B1 => n7823, B2 => n3186
                           , ZN => n1426);
   U563 : OAI22_X1 port map( A1 => n8480, A2 => n8800, B1 => n7824, B2 => n3186
                           , ZN => n1427);
   U564 : OAI22_X1 port map( A1 => n8480, A2 => n8803, B1 => n7825, B2 => n3186
                           , ZN => n1428);
   U565 : OAI22_X1 port map( A1 => n8480, A2 => n8806, B1 => n7826, B2 => n3186
                           , ZN => n1429);
   U566 : OAI22_X1 port map( A1 => n8481, A2 => n8809, B1 => n7827, B2 => n3186
                           , ZN => n1430);
   U567 : OAI22_X1 port map( A1 => n8481, A2 => n8821, B1 => n7828, B2 => n3186
                           , ZN => n1431);
   U568 : OAI22_X1 port map( A1 => n8497, A2 => n8791, B1 => n7901, B2 => n3184
                           , ZN => n1488);
   U569 : OAI22_X1 port map( A1 => n8498, A2 => n8794, B1 => n7902, B2 => n3184
                           , ZN => n1489);
   U570 : OAI22_X1 port map( A1 => n8498, A2 => n8797, B1 => n7903, B2 => n3184
                           , ZN => n1490);
   U571 : OAI22_X1 port map( A1 => n8498, A2 => n8800, B1 => n7904, B2 => n3184
                           , ZN => n1491);
   U572 : OAI22_X1 port map( A1 => n8498, A2 => n8803, B1 => n7905, B2 => n3184
                           , ZN => n1492);
   U573 : OAI22_X1 port map( A1 => n8498, A2 => n8806, B1 => n7906, B2 => n3184
                           , ZN => n1493);
   U574 : OAI22_X1 port map( A1 => n8499, A2 => n8809, B1 => n7907, B2 => n3184
                           , ZN => n1494);
   U575 : OAI22_X1 port map( A1 => n8499, A2 => n8821, B1 => n7908, B2 => n3184
                           , ZN => n1495);
   U576 : OAI22_X1 port map( A1 => n8524, A2 => n8790, B1 => n7805, B2 => n3180
                           , ZN => n1584);
   U577 : OAI22_X1 port map( A1 => n8525, A2 => n8793, B1 => n7807, B2 => n3180
                           , ZN => n1585);
   U578 : OAI22_X1 port map( A1 => n8525, A2 => n8796, B1 => n7809, B2 => n3180
                           , ZN => n1586);
   U579 : OAI22_X1 port map( A1 => n8525, A2 => n8799, B1 => n7811, B2 => n3180
                           , ZN => n1587);
   U580 : OAI22_X1 port map( A1 => n8525, A2 => n8802, B1 => n7813, B2 => n3180
                           , ZN => n1588);
   U581 : OAI22_X1 port map( A1 => n8525, A2 => n8805, B1 => n7815, B2 => n3180
                           , ZN => n1589);
   U582 : OAI22_X1 port map( A1 => n8526, A2 => n8808, B1 => n7817, B2 => n3180
                           , ZN => n1590);
   U583 : OAI22_X1 port map( A1 => n8526, A2 => n8820, B1 => n7819, B2 => n3180
                           , ZN => n1591);
   U584 : OAI22_X1 port map( A1 => n8542, A2 => n8790, B1 => n7917, B2 => n3178
                           , ZN => n1648);
   U585 : OAI22_X1 port map( A1 => n8543, A2 => n8793, B1 => n7918, B2 => n3178
                           , ZN => n1649);
   U586 : OAI22_X1 port map( A1 => n8543, A2 => n8796, B1 => n7919, B2 => n3178
                           , ZN => n1650);
   U587 : OAI22_X1 port map( A1 => n8543, A2 => n8799, B1 => n7920, B2 => n3178
                           , ZN => n1651);
   U588 : OAI22_X1 port map( A1 => n8543, A2 => n8802, B1 => n7921, B2 => n3178
                           , ZN => n1652);
   U589 : OAI22_X1 port map( A1 => n8543, A2 => n8805, B1 => n7922, B2 => n3178
                           , ZN => n1653);
   U590 : OAI22_X1 port map( A1 => n8544, A2 => n8808, B1 => n7923, B2 => n3178
                           , ZN => n1654);
   U591 : OAI22_X1 port map( A1 => n8544, A2 => n8820, B1 => n7924, B2 => n3178
                           , ZN => n1655);
   U592 : OAI22_X1 port map( A1 => n8569, A2 => n8790, B1 => n7853, B2 => n3175
                           , ZN => n1744);
   U593 : OAI22_X1 port map( A1 => n8570, A2 => n8793, B1 => n7854, B2 => n3175
                           , ZN => n1745);
   U594 : OAI22_X1 port map( A1 => n8570, A2 => n8796, B1 => n7855, B2 => n3175
                           , ZN => n1746);
   U595 : OAI22_X1 port map( A1 => n8570, A2 => n8799, B1 => n7856, B2 => n3175
                           , ZN => n1747);
   U596 : OAI22_X1 port map( A1 => n8570, A2 => n8802, B1 => n7857, B2 => n3175
                           , ZN => n1748);
   U597 : OAI22_X1 port map( A1 => n8570, A2 => n8805, B1 => n7858, B2 => n3175
                           , ZN => n1749);
   U598 : OAI22_X1 port map( A1 => n8571, A2 => n8808, B1 => n7859, B2 => n3175
                           , ZN => n1750);
   U599 : OAI22_X1 port map( A1 => n8571, A2 => n8820, B1 => n7860, B2 => n3175
                           , ZN => n1751);
   U600 : OAI22_X1 port map( A1 => n8578, A2 => n8790, B1 => n7689, B2 => n3173
                           , ZN => n1776);
   U601 : OAI22_X1 port map( A1 => n8579, A2 => n8793, B1 => n7690, B2 => n3173
                           , ZN => n1777);
   U602 : OAI22_X1 port map( A1 => n8579, A2 => n8796, B1 => n7691, B2 => n3173
                           , ZN => n1778);
   U603 : OAI22_X1 port map( A1 => n8579, A2 => n8799, B1 => n7692, B2 => n3173
                           , ZN => n1779);
   U604 : OAI22_X1 port map( A1 => n8579, A2 => n8802, B1 => n7693, B2 => n3173
                           , ZN => n1780);
   U605 : OAI22_X1 port map( A1 => n8579, A2 => n8805, B1 => n7694, B2 => n3173
                           , ZN => n1781);
   U606 : OAI22_X1 port map( A1 => n8580, A2 => n8808, B1 => n7695, B2 => n3173
                           , ZN => n1782);
   U607 : OAI22_X1 port map( A1 => n8580, A2 => n8820, B1 => n7696, B2 => n3173
                           , ZN => n1783);
   U608 : OAI22_X1 port map( A1 => n8587, A2 => n8790, B1 => n7681, B2 => n3172
                           , ZN => n1808);
   U609 : OAI22_X1 port map( A1 => n8588, A2 => n8793, B1 => n7682, B2 => n3172
                           , ZN => n1809);
   U610 : OAI22_X1 port map( A1 => n8588, A2 => n8796, B1 => n7683, B2 => n3172
                           , ZN => n1810);
   U611 : OAI22_X1 port map( A1 => n8588, A2 => n8799, B1 => n7684, B2 => n3172
                           , ZN => n1811);
   U612 : OAI22_X1 port map( A1 => n8588, A2 => n8802, B1 => n7685, B2 => n3172
                           , ZN => n1812);
   U613 : OAI22_X1 port map( A1 => n8588, A2 => n8805, B1 => n7686, B2 => n3172
                           , ZN => n1813);
   U614 : OAI22_X1 port map( A1 => n8589, A2 => n8808, B1 => n7687, B2 => n3172
                           , ZN => n1814);
   U615 : OAI22_X1 port map( A1 => n8589, A2 => n8820, B1 => n7688, B2 => n3172
                           , ZN => n1815);
   U616 : OAI22_X1 port map( A1 => n8632, A2 => n8789, B1 => n7761, B2 => n3167
                           , ZN => n1968);
   U617 : OAI22_X1 port map( A1 => n8633, A2 => n8792, B1 => n7762, B2 => n3167
                           , ZN => n1969);
   U618 : OAI22_X1 port map( A1 => n8633, A2 => n8795, B1 => n7763, B2 => n3167
                           , ZN => n1970);
   U619 : OAI22_X1 port map( A1 => n8633, A2 => n8798, B1 => n7764, B2 => n3167
                           , ZN => n1971);
   U620 : OAI22_X1 port map( A1 => n8633, A2 => n8801, B1 => n7765, B2 => n3167
                           , ZN => n1972);
   U621 : OAI22_X1 port map( A1 => n8633, A2 => n8804, B1 => n7766, B2 => n3167
                           , ZN => n1973);
   U622 : OAI22_X1 port map( A1 => n8634, A2 => n8807, B1 => n7767, B2 => n3167
                           , ZN => n1974);
   U623 : OAI22_X1 port map( A1 => n8634, A2 => n8819, B1 => n7768, B2 => n3167
                           , ZN => n1975);
   U624 : OAI22_X1 port map( A1 => n8650, A2 => n8789, B1 => n7697, B2 => n3164
                           , ZN => n2032);
   U625 : OAI22_X1 port map( A1 => n8651, A2 => n8792, B1 => n7698, B2 => n3164
                           , ZN => n2033);
   U626 : OAI22_X1 port map( A1 => n8651, A2 => n8795, B1 => n7699, B2 => n3164
                           , ZN => n2034);
   U627 : OAI22_X1 port map( A1 => n8651, A2 => n8798, B1 => n7700, B2 => n3164
                           , ZN => n2035);
   U628 : OAI22_X1 port map( A1 => n8651, A2 => n8801, B1 => n7701, B2 => n3164
                           , ZN => n2036);
   U629 : OAI22_X1 port map( A1 => n8651, A2 => n8804, B1 => n7702, B2 => n3164
                           , ZN => n2037);
   U630 : OAI22_X1 port map( A1 => n8652, A2 => n8807, B1 => n7703, B2 => n3164
                           , ZN => n2038);
   U631 : OAI22_X1 port map( A1 => n8652, A2 => n8819, B1 => n7704, B2 => n3164
                           , ZN => n2039);
   U632 : OAI22_X1 port map( A1 => n8659, A2 => n8789, B1 => n7806, B2 => n3162
                           , ZN => n2064);
   U633 : OAI22_X1 port map( A1 => n8660, A2 => n8792, B1 => n7808, B2 => n3162
                           , ZN => n2065);
   U634 : OAI22_X1 port map( A1 => n8660, A2 => n8795, B1 => n7810, B2 => n3162
                           , ZN => n2066);
   U635 : OAI22_X1 port map( A1 => n8660, A2 => n8798, B1 => n7812, B2 => n3162
                           , ZN => n2067);
   U636 : OAI22_X1 port map( A1 => n8660, A2 => n8801, B1 => n7814, B2 => n3162
                           , ZN => n2068);
   U637 : OAI22_X1 port map( A1 => n8660, A2 => n8804, B1 => n7816, B2 => n3162
                           , ZN => n2069);
   U638 : OAI22_X1 port map( A1 => n8661, A2 => n8807, B1 => n7818, B2 => n3162
                           , ZN => n2070);
   U639 : OAI22_X1 port map( A1 => n8661, A2 => n8819, B1 => n7820, B2 => n3162
                           , ZN => n2071);
   U640 : OAI22_X1 port map( A1 => n8668, A2 => n8789, B1 => n7869, B2 => n3160
                           , ZN => n2096);
   U641 : OAI22_X1 port map( A1 => n8669, A2 => n8792, B1 => n7870, B2 => n3160
                           , ZN => n2097);
   U642 : OAI22_X1 port map( A1 => n8669, A2 => n8795, B1 => n7871, B2 => n3160
                           , ZN => n2098);
   U643 : OAI22_X1 port map( A1 => n8669, A2 => n8798, B1 => n7872, B2 => n3160
                           , ZN => n2099);
   U644 : OAI22_X1 port map( A1 => n8669, A2 => n8801, B1 => n7873, B2 => n3160
                           , ZN => n2100);
   U645 : OAI22_X1 port map( A1 => n8669, A2 => n8804, B1 => n7874, B2 => n3160
                           , ZN => n2101);
   U646 : OAI22_X1 port map( A1 => n8670, A2 => n8807, B1 => n7875, B2 => n3160
                           , ZN => n2102);
   U647 : OAI22_X1 port map( A1 => n8670, A2 => n8819, B1 => n7876, B2 => n3160
                           , ZN => n2103);
   U648 : OAI22_X1 port map( A1 => n8695, A2 => n8789, B1 => n7753, B2 => n3154
                           , ZN => n2192);
   U649 : OAI22_X1 port map( A1 => n8696, A2 => n8792, B1 => n7754, B2 => n3154
                           , ZN => n2193);
   U650 : OAI22_X1 port map( A1 => n8696, A2 => n8795, B1 => n7755, B2 => n3154
                           , ZN => n2194);
   U651 : OAI22_X1 port map( A1 => n8696, A2 => n8798, B1 => n7756, B2 => n3154
                           , ZN => n2195);
   U652 : OAI22_X1 port map( A1 => n8696, A2 => n8801, B1 => n7757, B2 => n3154
                           , ZN => n2196);
   U653 : OAI22_X1 port map( A1 => n8696, A2 => n8804, B1 => n7758, B2 => n3154
                           , ZN => n2197);
   U654 : OAI22_X1 port map( A1 => n8697, A2 => n8807, B1 => n7759, B2 => n3154
                           , ZN => n2198);
   U655 : OAI22_X1 port map( A1 => n8697, A2 => n8819, B1 => n7760, B2 => n3154
                           , ZN => n2199);
   U656 : OAI22_X1 port map( A1 => n8704, A2 => n8789, B1 => n7637, B2 => n3152
                           , ZN => n2224);
   U657 : OAI22_X1 port map( A1 => n8705, A2 => n8792, B1 => n7638, B2 => n3152
                           , ZN => n2225);
   U658 : OAI22_X1 port map( A1 => n8705, A2 => n8795, B1 => n7639, B2 => n3152
                           , ZN => n2226);
   U659 : OAI22_X1 port map( A1 => n8705, A2 => n8798, B1 => n7640, B2 => n3152
                           , ZN => n2227);
   U660 : OAI22_X1 port map( A1 => n8705, A2 => n8801, B1 => n7641, B2 => n3152
                           , ZN => n2228);
   U661 : OAI22_X1 port map( A1 => n8705, A2 => n8804, B1 => n7642, B2 => n3152
                           , ZN => n2229);
   U662 : OAI22_X1 port map( A1 => n8706, A2 => n8807, B1 => n7643, B2 => n3152
                           , ZN => n2230);
   U663 : OAI22_X1 port map( A1 => n8706, A2 => n8819, B1 => n7644, B2 => n3152
                           , ZN => n2231);
   U664 : OAI22_X1 port map( A1 => n8713, A2 => n8789, B1 => n7861, B2 => n3150
                           , ZN => n2256);
   U665 : OAI22_X1 port map( A1 => n8714, A2 => n8792, B1 => n7862, B2 => n3150
                           , ZN => n2257);
   U666 : OAI22_X1 port map( A1 => n8714, A2 => n8795, B1 => n7863, B2 => n3150
                           , ZN => n2258);
   U667 : OAI22_X1 port map( A1 => n8714, A2 => n8798, B1 => n7864, B2 => n3150
                           , ZN => n2259);
   U668 : OAI22_X1 port map( A1 => n8714, A2 => n8801, B1 => n7865, B2 => n3150
                           , ZN => n2260);
   U669 : OAI22_X1 port map( A1 => n8714, A2 => n8804, B1 => n7866, B2 => n3150
                           , ZN => n2261);
   U670 : OAI22_X1 port map( A1 => n8715, A2 => n8807, B1 => n7867, B2 => n3150
                           , ZN => n2262);
   U671 : OAI22_X1 port map( A1 => n8715, A2 => n8819, B1 => n7868, B2 => n3150
                           , ZN => n2263);
   U672 : OAI22_X1 port map( A1 => n8815, A2 => n8789, B1 => n7909, B2 => n3116
                           , ZN => n2288);
   U673 : OAI22_X1 port map( A1 => n8816, A2 => n8792, B1 => n7910, B2 => n3116
                           , ZN => n2289);
   U674 : OAI22_X1 port map( A1 => n8816, A2 => n8795, B1 => n7911, B2 => n3116
                           , ZN => n2290);
   U675 : OAI22_X1 port map( A1 => n8816, A2 => n8798, B1 => n7912, B2 => n3116
                           , ZN => n2291);
   U676 : OAI22_X1 port map( A1 => n8816, A2 => n8801, B1 => n7913, B2 => n3116
                           , ZN => n2292);
   U677 : OAI22_X1 port map( A1 => n8816, A2 => n8804, B1 => n7914, B2 => n3116
                           , ZN => n2293);
   U678 : OAI22_X1 port map( A1 => n8817, A2 => n8807, B1 => n7915, B2 => n3116
                           , ZN => n2294);
   U679 : OAI22_X1 port map( A1 => n8817, A2 => n8819, B1 => n7916, B2 => n3116
                           , ZN => n2295);
   U680 : OAI22_X1 port map( A1 => n7997, A2 => n3190, B1 => n8438, B2 => n8719
                           , ZN => n1272);
   U681 : OAI22_X1 port map( A1 => n7998, A2 => n8437, B1 => n8438, B2 => n8722
                           , ZN => n1273);
   U682 : OAI22_X1 port map( A1 => n7999, A2 => n8437, B1 => n8438, B2 => n8725
                           , ZN => n1274);
   U683 : OAI22_X1 port map( A1 => n8000, A2 => n8437, B1 => n8438, B2 => n8728
                           , ZN => n1275);
   U684 : OAI22_X1 port map( A1 => n8001, A2 => n8437, B1 => n8439, B2 => n8731
                           , ZN => n1276);
   U685 : OAI22_X1 port map( A1 => n8002, A2 => n8437, B1 => n8439, B2 => n8734
                           , ZN => n1277);
   U686 : OAI22_X1 port map( A1 => n8003, A2 => n8437, B1 => n8439, B2 => n8737
                           , ZN => n1278);
   U687 : OAI22_X1 port map( A1 => n8004, A2 => n8437, B1 => n8439, B2 => n8740
                           , ZN => n1279);
   U688 : OAI22_X1 port map( A1 => n8005, A2 => n8437, B1 => n8440, B2 => n8743
                           , ZN => n1280);
   U689 : OAI22_X1 port map( A1 => n8006, A2 => n8437, B1 => n8440, B2 => n8746
                           , ZN => n1281);
   U690 : OAI22_X1 port map( A1 => n8007, A2 => n8437, B1 => n8440, B2 => n8749
                           , ZN => n1282);
   U691 : OAI22_X1 port map( A1 => n8008, A2 => n8437, B1 => n8440, B2 => n8752
                           , ZN => n1283);
   U692 : OAI22_X1 port map( A1 => n8009, A2 => n3190, B1 => n8441, B2 => n8755
                           , ZN => n1284);
   U693 : OAI22_X1 port map( A1 => n8010, A2 => n8437, B1 => n8441, B2 => n8758
                           , ZN => n1285);
   U694 : OAI22_X1 port map( A1 => n8011, A2 => n3190, B1 => n8441, B2 => n8761
                           , ZN => n1286);
   U695 : OAI22_X1 port map( A1 => n8012, A2 => n8437, B1 => n8441, B2 => n8764
                           , ZN => n1287);
   U696 : OAI22_X1 port map( A1 => n8013, A2 => n3190, B1 => n8442, B2 => n8767
                           , ZN => n1288);
   U697 : OAI22_X1 port map( A1 => n8014, A2 => n8437, B1 => n8442, B2 => n8770
                           , ZN => n1289);
   U698 : OAI22_X1 port map( A1 => n8015, A2 => n3190, B1 => n8442, B2 => n8773
                           , ZN => n1290);
   U699 : OAI22_X1 port map( A1 => n8016, A2 => n8437, B1 => n8442, B2 => n8776
                           , ZN => n1291);
   U700 : OAI22_X1 port map( A1 => n8017, A2 => n3190, B1 => n8443, B2 => n8779
                           , ZN => n1292);
   U701 : OAI22_X1 port map( A1 => n8018, A2 => n8437, B1 => n8443, B2 => n8782
                           , ZN => n1293);
   U702 : OAI22_X1 port map( A1 => n8019, A2 => n3190, B1 => n8443, B2 => n8785
                           , ZN => n1294);
   U703 : OAI22_X1 port map( A1 => n8020, A2 => n8437, B1 => n8443, B2 => n8788
                           , ZN => n1295);
   U704 : OAI22_X1 port map( A1 => n8021, A2 => n3190, B1 => n8444, B2 => n8791
                           , ZN => n1296);
   U705 : OAI22_X1 port map( A1 => n8022, A2 => n8437, B1 => n8444, B2 => n8794
                           , ZN => n1297);
   U706 : OAI22_X1 port map( A1 => n8023, A2 => n3190, B1 => n8444, B2 => n8797
                           , ZN => n1298);
   U707 : OAI22_X1 port map( A1 => n8024, A2 => n8437, B1 => n8444, B2 => n8800
                           , ZN => n1299);
   U708 : OAI22_X1 port map( A1 => n8025, A2 => n3190, B1 => n8445, B2 => n8803
                           , ZN => n1300);
   U709 : OAI22_X1 port map( A1 => n8026, A2 => n8437, B1 => n8445, B2 => n8806
                           , ZN => n1301);
   U710 : OAI22_X1 port map( A1 => n8027, A2 => n3190, B1 => n8445, B2 => n8809
                           , ZN => n1302);
   U711 : OAI22_X1 port map( A1 => n8028, A2 => n8437, B1 => n8445, B2 => n8821
                           , ZN => n1303);
   U712 : OAI22_X1 port map( A1 => n8475, A2 => n8719, B1 => n8029, B2 => n8474
                           , ZN => n1400);
   U713 : OAI22_X1 port map( A1 => n8475, A2 => n8722, B1 => n8030, B2 => n8474
                           , ZN => n1401);
   U714 : OAI22_X1 port map( A1 => n8475, A2 => n8725, B1 => n8031, B2 => n8474
                           , ZN => n1402);
   U715 : OAI22_X1 port map( A1 => n8475, A2 => n8728, B1 => n8032, B2 => n8474
                           , ZN => n1403);
   U716 : OAI22_X1 port map( A1 => n8475, A2 => n8731, B1 => n8033, B2 => n8474
                           , ZN => n1404);
   U717 : OAI22_X1 port map( A1 => n8476, A2 => n8734, B1 => n8034, B2 => n8474
                           , ZN => n1405);
   U718 : OAI22_X1 port map( A1 => n8476, A2 => n8737, B1 => n8035, B2 => n8474
                           , ZN => n1406);
   U719 : OAI22_X1 port map( A1 => n8476, A2 => n8740, B1 => n8036, B2 => n8474
                           , ZN => n1407);
   U720 : OAI22_X1 port map( A1 => n8476, A2 => n8743, B1 => n8037, B2 => n8474
                           , ZN => n1408);
   U721 : OAI22_X1 port map( A1 => n8476, A2 => n8746, B1 => n8038, B2 => n8474
                           , ZN => n1409);
   U722 : OAI22_X1 port map( A1 => n8477, A2 => n8749, B1 => n8039, B2 => n8474
                           , ZN => n1410);
   U723 : OAI22_X1 port map( A1 => n8477, A2 => n8752, B1 => n8040, B2 => n8474
                           , ZN => n1411);
   U724 : OAI22_X1 port map( A1 => n8477, A2 => n8755, B1 => n8041, B2 => n3186
                           , ZN => n1412);
   U725 : OAI22_X1 port map( A1 => n8477, A2 => n8758, B1 => n8042, B2 => n3186
                           , ZN => n1413);
   U726 : OAI22_X1 port map( A1 => n8477, A2 => n8761, B1 => n8043, B2 => n3186
                           , ZN => n1414);
   U727 : OAI22_X1 port map( A1 => n8478, A2 => n8764, B1 => n8044, B2 => n8474
                           , ZN => n1415);
   U728 : OAI22_X1 port map( A1 => n8478, A2 => n8767, B1 => n8045, B2 => n8474
                           , ZN => n1416);
   U729 : OAI22_X1 port map( A1 => n8478, A2 => n8770, B1 => n8046, B2 => n8474
                           , ZN => n1417);
   U730 : OAI22_X1 port map( A1 => n8478, A2 => n8773, B1 => n8047, B2 => n8474
                           , ZN => n1418);
   U731 : OAI22_X1 port map( A1 => n8478, A2 => n8776, B1 => n8048, B2 => n8474
                           , ZN => n1419);
   U732 : OAI22_X1 port map( A1 => n8479, A2 => n8779, B1 => n8049, B2 => n8474
                           , ZN => n1420);
   U733 : OAI22_X1 port map( A1 => n8479, A2 => n8782, B1 => n8050, B2 => n8474
                           , ZN => n1421);
   U734 : OAI22_X1 port map( A1 => n8479, A2 => n8785, B1 => n8051, B2 => n8474
                           , ZN => n1422);
   U735 : OAI22_X1 port map( A1 => n8479, A2 => n8788, B1 => n8052, B2 => n8474
                           , ZN => n1423);
   U736 : OAI22_X1 port map( A1 => n8493, A2 => n8719, B1 => n8157, B2 => n8492
                           , ZN => n1464);
   U737 : OAI22_X1 port map( A1 => n8493, A2 => n8722, B1 => n8158, B2 => n8492
                           , ZN => n1465);
   U738 : OAI22_X1 port map( A1 => n8493, A2 => n8725, B1 => n8159, B2 => n8492
                           , ZN => n1466);
   U739 : OAI22_X1 port map( A1 => n8493, A2 => n8728, B1 => n8160, B2 => n8492
                           , ZN => n1467);
   U740 : OAI22_X1 port map( A1 => n8493, A2 => n8731, B1 => n8161, B2 => n8492
                           , ZN => n1468);
   U741 : OAI22_X1 port map( A1 => n8494, A2 => n8734, B1 => n8162, B2 => n8492
                           , ZN => n1469);
   U742 : OAI22_X1 port map( A1 => n8494, A2 => n8737, B1 => n8163, B2 => n8492
                           , ZN => n1470);
   U743 : OAI22_X1 port map( A1 => n8494, A2 => n8740, B1 => n8164, B2 => n8492
                           , ZN => n1471);
   U744 : OAI22_X1 port map( A1 => n8494, A2 => n8743, B1 => n8165, B2 => n8492
                           , ZN => n1472);
   U745 : OAI22_X1 port map( A1 => n8494, A2 => n8746, B1 => n8166, B2 => n8492
                           , ZN => n1473);
   U746 : OAI22_X1 port map( A1 => n8495, A2 => n8749, B1 => n8167, B2 => n8492
                           , ZN => n1474);
   U747 : OAI22_X1 port map( A1 => n8495, A2 => n8752, B1 => n8168, B2 => n8492
                           , ZN => n1475);
   U748 : OAI22_X1 port map( A1 => n8495, A2 => n8755, B1 => n8169, B2 => n3184
                           , ZN => n1476);
   U749 : OAI22_X1 port map( A1 => n8495, A2 => n8758, B1 => n8170, B2 => n3184
                           , ZN => n1477);
   U750 : OAI22_X1 port map( A1 => n8495, A2 => n8761, B1 => n8171, B2 => n3184
                           , ZN => n1478);
   U751 : OAI22_X1 port map( A1 => n8496, A2 => n8764, B1 => n8172, B2 => n8492
                           , ZN => n1479);
   U752 : OAI22_X1 port map( A1 => n8496, A2 => n8767, B1 => n8173, B2 => n8492
                           , ZN => n1480);
   U753 : OAI22_X1 port map( A1 => n8496, A2 => n8770, B1 => n8174, B2 => n8492
                           , ZN => n1481);
   U754 : OAI22_X1 port map( A1 => n8496, A2 => n8773, B1 => n8175, B2 => n8492
                           , ZN => n1482);
   U755 : OAI22_X1 port map( A1 => n8496, A2 => n8776, B1 => n8176, B2 => n8492
                           , ZN => n1483);
   U756 : OAI22_X1 port map( A1 => n8497, A2 => n8779, B1 => n8177, B2 => n8492
                           , ZN => n1484);
   U757 : OAI22_X1 port map( A1 => n8497, A2 => n8782, B1 => n8178, B2 => n8492
                           , ZN => n1485);
   U758 : OAI22_X1 port map( A1 => n8497, A2 => n8785, B1 => n8179, B2 => n8492
                           , ZN => n1486);
   U759 : OAI22_X1 port map( A1 => n8497, A2 => n8788, B1 => n8180, B2 => n8492
                           , ZN => n1487);
   U760 : OAI22_X1 port map( A1 => n8520, A2 => n8718, B1 => n7973, B2 => n8519
                           , ZN => n1560);
   U761 : OAI22_X1 port map( A1 => n8520, A2 => n8721, B1 => n7974, B2 => n8519
                           , ZN => n1561);
   U762 : OAI22_X1 port map( A1 => n8520, A2 => n8724, B1 => n7975, B2 => n8519
                           , ZN => n1562);
   U763 : OAI22_X1 port map( A1 => n8520, A2 => n8727, B1 => n7976, B2 => n8519
                           , ZN => n1563);
   U764 : OAI22_X1 port map( A1 => n8520, A2 => n8730, B1 => n7977, B2 => n8519
                           , ZN => n1564);
   U765 : OAI22_X1 port map( A1 => n8521, A2 => n8733, B1 => n7978, B2 => n8519
                           , ZN => n1565);
   U766 : OAI22_X1 port map( A1 => n8521, A2 => n8736, B1 => n7979, B2 => n8519
                           , ZN => n1566);
   U767 : OAI22_X1 port map( A1 => n8521, A2 => n8739, B1 => n7980, B2 => n8519
                           , ZN => n1567);
   U768 : OAI22_X1 port map( A1 => n8521, A2 => n8742, B1 => n7981, B2 => n8519
                           , ZN => n1568);
   U769 : OAI22_X1 port map( A1 => n8521, A2 => n8745, B1 => n7982, B2 => n8519
                           , ZN => n1569);
   U770 : OAI22_X1 port map( A1 => n8522, A2 => n8748, B1 => n7983, B2 => n8519
                           , ZN => n1570);
   U771 : OAI22_X1 port map( A1 => n8522, A2 => n8751, B1 => n7984, B2 => n8519
                           , ZN => n1571);
   U772 : OAI22_X1 port map( A1 => n8522, A2 => n8754, B1 => n7985, B2 => n3180
                           , ZN => n1572);
   U773 : OAI22_X1 port map( A1 => n8522, A2 => n8757, B1 => n7986, B2 => n3180
                           , ZN => n1573);
   U774 : OAI22_X1 port map( A1 => n8522, A2 => n8760, B1 => n7987, B2 => n3180
                           , ZN => n1574);
   U775 : OAI22_X1 port map( A1 => n8523, A2 => n8763, B1 => n7988, B2 => n8519
                           , ZN => n1575);
   U776 : OAI22_X1 port map( A1 => n8523, A2 => n8766, B1 => n7989, B2 => n8519
                           , ZN => n1576);
   U777 : OAI22_X1 port map( A1 => n8523, A2 => n8769, B1 => n7990, B2 => n8519
                           , ZN => n1577);
   U778 : OAI22_X1 port map( A1 => n8523, A2 => n8772, B1 => n7991, B2 => n8519
                           , ZN => n1578);
   U779 : OAI22_X1 port map( A1 => n8523, A2 => n8775, B1 => n7992, B2 => n8519
                           , ZN => n1579);
   U780 : OAI22_X1 port map( A1 => n8524, A2 => n8778, B1 => n7993, B2 => n8519
                           , ZN => n1580);
   U781 : OAI22_X1 port map( A1 => n8524, A2 => n8781, B1 => n7994, B2 => n8519
                           , ZN => n1581);
   U782 : OAI22_X1 port map( A1 => n8524, A2 => n8784, B1 => n7995, B2 => n8519
                           , ZN => n1582);
   U783 : OAI22_X1 port map( A1 => n8524, A2 => n8787, B1 => n7996, B2 => n8519
                           , ZN => n1583);
   U784 : OAI22_X1 port map( A1 => n8538, A2 => n8718, B1 => n8205, B2 => n8537
                           , ZN => n1624);
   U785 : OAI22_X1 port map( A1 => n8538, A2 => n8721, B1 => n8206, B2 => n8537
                           , ZN => n1625);
   U786 : OAI22_X1 port map( A1 => n8538, A2 => n8724, B1 => n8207, B2 => n8537
                           , ZN => n1626);
   U787 : OAI22_X1 port map( A1 => n8538, A2 => n8727, B1 => n8208, B2 => n8537
                           , ZN => n1627);
   U788 : OAI22_X1 port map( A1 => n8538, A2 => n8730, B1 => n8209, B2 => n8537
                           , ZN => n1628);
   U789 : OAI22_X1 port map( A1 => n8539, A2 => n8733, B1 => n8210, B2 => n8537
                           , ZN => n1629);
   U790 : OAI22_X1 port map( A1 => n8539, A2 => n8736, B1 => n8211, B2 => n8537
                           , ZN => n1630);
   U791 : OAI22_X1 port map( A1 => n8539, A2 => n8739, B1 => n8212, B2 => n8537
                           , ZN => n1631);
   U792 : OAI22_X1 port map( A1 => n8539, A2 => n8742, B1 => n8213, B2 => n8537
                           , ZN => n1632);
   U793 : OAI22_X1 port map( A1 => n8539, A2 => n8745, B1 => n8214, B2 => n8537
                           , ZN => n1633);
   U794 : OAI22_X1 port map( A1 => n8540, A2 => n8748, B1 => n8215, B2 => n8537
                           , ZN => n1634);
   U795 : OAI22_X1 port map( A1 => n8540, A2 => n8751, B1 => n8216, B2 => n8537
                           , ZN => n1635);
   U796 : OAI22_X1 port map( A1 => n8540, A2 => n8754, B1 => n8217, B2 => n3178
                           , ZN => n1636);
   U797 : OAI22_X1 port map( A1 => n8540, A2 => n8757, B1 => n8218, B2 => n3178
                           , ZN => n1637);
   U798 : OAI22_X1 port map( A1 => n8540, A2 => n8760, B1 => n8219, B2 => n3178
                           , ZN => n1638);
   U799 : OAI22_X1 port map( A1 => n8541, A2 => n8763, B1 => n8220, B2 => n8537
                           , ZN => n1639);
   U800 : OAI22_X1 port map( A1 => n8541, A2 => n8766, B1 => n8221, B2 => n8537
                           , ZN => n1640);
   U801 : OAI22_X1 port map( A1 => n8541, A2 => n8769, B1 => n8222, B2 => n8537
                           , ZN => n1641);
   U802 : OAI22_X1 port map( A1 => n8541, A2 => n8772, B1 => n8223, B2 => n8537
                           , ZN => n1642);
   U803 : OAI22_X1 port map( A1 => n8541, A2 => n8775, B1 => n8224, B2 => n8537
                           , ZN => n1643);
   U804 : OAI22_X1 port map( A1 => n8542, A2 => n8778, B1 => n8225, B2 => n8537
                           , ZN => n1644);
   U805 : OAI22_X1 port map( A1 => n8542, A2 => n8781, B1 => n8226, B2 => n8537
                           , ZN => n1645);
   U806 : OAI22_X1 port map( A1 => n8542, A2 => n8784, B1 => n8227, B2 => n8537
                           , ZN => n1646);
   U807 : OAI22_X1 port map( A1 => n8542, A2 => n8787, B1 => n8228, B2 => n8537
                           , ZN => n1647);
   U808 : OAI22_X1 port map( A1 => n8565, A2 => n8718, B1 => n8085, B2 => n8564
                           , ZN => n1720);
   U809 : OAI22_X1 port map( A1 => n8565, A2 => n8721, B1 => n8086, B2 => n8564
                           , ZN => n1721);
   U810 : OAI22_X1 port map( A1 => n8565, A2 => n8724, B1 => n8087, B2 => n8564
                           , ZN => n1722);
   U811 : OAI22_X1 port map( A1 => n8565, A2 => n8727, B1 => n8088, B2 => n8564
                           , ZN => n1723);
   U812 : OAI22_X1 port map( A1 => n8565, A2 => n8730, B1 => n8089, B2 => n8564
                           , ZN => n1724);
   U813 : OAI22_X1 port map( A1 => n8566, A2 => n8733, B1 => n8090, B2 => n8564
                           , ZN => n1725);
   U814 : OAI22_X1 port map( A1 => n8566, A2 => n8736, B1 => n8091, B2 => n8564
                           , ZN => n1726);
   U815 : OAI22_X1 port map( A1 => n8566, A2 => n8739, B1 => n8092, B2 => n8564
                           , ZN => n1727);
   U816 : OAI22_X1 port map( A1 => n8566, A2 => n8742, B1 => n8093, B2 => n8564
                           , ZN => n1728);
   U817 : OAI22_X1 port map( A1 => n8566, A2 => n8745, B1 => n8094, B2 => n8564
                           , ZN => n1729);
   U818 : OAI22_X1 port map( A1 => n8567, A2 => n8748, B1 => n8095, B2 => n8564
                           , ZN => n1730);
   U819 : OAI22_X1 port map( A1 => n8567, A2 => n8751, B1 => n8096, B2 => n8564
                           , ZN => n1731);
   U820 : OAI22_X1 port map( A1 => n8567, A2 => n8754, B1 => n8097, B2 => n3175
                           , ZN => n1732);
   U821 : OAI22_X1 port map( A1 => n8567, A2 => n8757, B1 => n8098, B2 => n3175
                           , ZN => n1733);
   U822 : OAI22_X1 port map( A1 => n8567, A2 => n8760, B1 => n8099, B2 => n3175
                           , ZN => n1734);
   U823 : OAI22_X1 port map( A1 => n8568, A2 => n8763, B1 => n8100, B2 => n8564
                           , ZN => n1735);
   U824 : OAI22_X1 port map( A1 => n8568, A2 => n8766, B1 => n8101, B2 => n8564
                           , ZN => n1736);
   U825 : OAI22_X1 port map( A1 => n8568, A2 => n8769, B1 => n8102, B2 => n8564
                           , ZN => n1737);
   U826 : OAI22_X1 port map( A1 => n8568, A2 => n8772, B1 => n8103, B2 => n8564
                           , ZN => n1738);
   U827 : OAI22_X1 port map( A1 => n8568, A2 => n8775, B1 => n8104, B2 => n8564
                           , ZN => n1739);
   U828 : OAI22_X1 port map( A1 => n8569, A2 => n8778, B1 => n8105, B2 => n8564
                           , ZN => n1740);
   U829 : OAI22_X1 port map( A1 => n8569, A2 => n8781, B1 => n8106, B2 => n8564
                           , ZN => n1741);
   U830 : OAI22_X1 port map( A1 => n8569, A2 => n8784, B1 => n8107, B2 => n8564
                           , ZN => n1742);
   U831 : OAI22_X1 port map( A1 => n8569, A2 => n8787, B1 => n8108, B2 => n8564
                           , ZN => n1743);
   U832 : OAI22_X1 port map( A1 => n8574, A2 => n8718, B1 => n7829, B2 => n8573
                           , ZN => n1752);
   U833 : OAI22_X1 port map( A1 => n8574, A2 => n8721, B1 => n7830, B2 => n8573
                           , ZN => n1753);
   U834 : OAI22_X1 port map( A1 => n8574, A2 => n8724, B1 => n7831, B2 => n8573
                           , ZN => n1754);
   U835 : OAI22_X1 port map( A1 => n8574, A2 => n8727, B1 => n7832, B2 => n8573
                           , ZN => n1755);
   U836 : OAI22_X1 port map( A1 => n8574, A2 => n8730, B1 => n7833, B2 => n8573
                           , ZN => n1756);
   U837 : OAI22_X1 port map( A1 => n8575, A2 => n8733, B1 => n7834, B2 => n8573
                           , ZN => n1757);
   U838 : OAI22_X1 port map( A1 => n8575, A2 => n8736, B1 => n7835, B2 => n8573
                           , ZN => n1758);
   U839 : OAI22_X1 port map( A1 => n8575, A2 => n8739, B1 => n7836, B2 => n8573
                           , ZN => n1759);
   U840 : OAI22_X1 port map( A1 => n8575, A2 => n8742, B1 => n7837, B2 => n8573
                           , ZN => n1760);
   U841 : OAI22_X1 port map( A1 => n8575, A2 => n8745, B1 => n7838, B2 => n8573
                           , ZN => n1761);
   U842 : OAI22_X1 port map( A1 => n8576, A2 => n8748, B1 => n7839, B2 => n8573
                           , ZN => n1762);
   U843 : OAI22_X1 port map( A1 => n8576, A2 => n8751, B1 => n7840, B2 => n8573
                           , ZN => n1763);
   U844 : OAI22_X1 port map( A1 => n8576, A2 => n8754, B1 => n7705, B2 => n3173
                           , ZN => n1764);
   U845 : OAI22_X1 port map( A1 => n8576, A2 => n8757, B1 => n7706, B2 => n3173
                           , ZN => n1765);
   U846 : OAI22_X1 port map( A1 => n8576, A2 => n8760, B1 => n7707, B2 => n3173
                           , ZN => n1766);
   U847 : OAI22_X1 port map( A1 => n8577, A2 => n8763, B1 => n7708, B2 => n8573
                           , ZN => n1767);
   U848 : OAI22_X1 port map( A1 => n8577, A2 => n8766, B1 => n7709, B2 => n8573
                           , ZN => n1768);
   U849 : OAI22_X1 port map( A1 => n8577, A2 => n8769, B1 => n7710, B2 => n8573
                           , ZN => n1769);
   U850 : OAI22_X1 port map( A1 => n8577, A2 => n8772, B1 => n7711, B2 => n8573
                           , ZN => n1770);
   U851 : OAI22_X1 port map( A1 => n8577, A2 => n8775, B1 => n7712, B2 => n8573
                           , ZN => n1771);
   U852 : OAI22_X1 port map( A1 => n8578, A2 => n8778, B1 => n7713, B2 => n8573
                           , ZN => n1772);
   U853 : OAI22_X1 port map( A1 => n8578, A2 => n8781, B1 => n7714, B2 => n8573
                           , ZN => n1773);
   U854 : OAI22_X1 port map( A1 => n8578, A2 => n8784, B1 => n7715, B2 => n8573
                           , ZN => n1774);
   U855 : OAI22_X1 port map( A1 => n8578, A2 => n8787, B1 => n7716, B2 => n8573
                           , ZN => n1775);
   U856 : OAI22_X1 port map( A1 => n8583, A2 => n8718, B1 => n7781, B2 => n8582
                           , ZN => n1784);
   U857 : OAI22_X1 port map( A1 => n8583, A2 => n8721, B1 => n7782, B2 => n8582
                           , ZN => n1785);
   U858 : OAI22_X1 port map( A1 => n8583, A2 => n8724, B1 => n7783, B2 => n8582
                           , ZN => n1786);
   U859 : OAI22_X1 port map( A1 => n8583, A2 => n8727, B1 => n7784, B2 => n8582
                           , ZN => n1787);
   U860 : OAI22_X1 port map( A1 => n8583, A2 => n8730, B1 => n7785, B2 => n8582
                           , ZN => n1788);
   U861 : OAI22_X1 port map( A1 => n8584, A2 => n8733, B1 => n7786, B2 => n8582
                           , ZN => n1789);
   U862 : OAI22_X1 port map( A1 => n8584, A2 => n8736, B1 => n7787, B2 => n8582
                           , ZN => n1790);
   U863 : OAI22_X1 port map( A1 => n8584, A2 => n8739, B1 => n7788, B2 => n8582
                           , ZN => n1791);
   U864 : OAI22_X1 port map( A1 => n8584, A2 => n8742, B1 => n7798, B2 => n8582
                           , ZN => n1792);
   U865 : OAI22_X1 port map( A1 => n8584, A2 => n8745, B1 => n7800, B2 => n8582
                           , ZN => n1793);
   U866 : OAI22_X1 port map( A1 => n8585, A2 => n8748, B1 => n7802, B2 => n8582
                           , ZN => n1794);
   U867 : OAI22_X1 port map( A1 => n8585, A2 => n8751, B1 => n7804, B2 => n8582
                           , ZN => n1795);
   U868 : OAI22_X1 port map( A1 => n8585, A2 => n8754, B1 => n7658, B2 => n3172
                           , ZN => n1796);
   U869 : OAI22_X1 port map( A1 => n8585, A2 => n8757, B1 => n7660, B2 => n3172
                           , ZN => n1797);
   U870 : OAI22_X1 port map( A1 => n8585, A2 => n8760, B1 => n7662, B2 => n3172
                           , ZN => n1798);
   U871 : OAI22_X1 port map( A1 => n8586, A2 => n8763, B1 => n7664, B2 => n8582
                           , ZN => n1799);
   U872 : OAI22_X1 port map( A1 => n8586, A2 => n8766, B1 => n7666, B2 => n8582
                           , ZN => n1800);
   U873 : OAI22_X1 port map( A1 => n8586, A2 => n8769, B1 => n7668, B2 => n8582
                           , ZN => n1801);
   U874 : OAI22_X1 port map( A1 => n8586, A2 => n8772, B1 => n7670, B2 => n8582
                           , ZN => n1802);
   U875 : OAI22_X1 port map( A1 => n8586, A2 => n8775, B1 => n7672, B2 => n8582
                           , ZN => n1803);
   U876 : OAI22_X1 port map( A1 => n8587, A2 => n8778, B1 => n7674, B2 => n8582
                           , ZN => n1804);
   U877 : OAI22_X1 port map( A1 => n8587, A2 => n8781, B1 => n7676, B2 => n8582
                           , ZN => n1805);
   U878 : OAI22_X1 port map( A1 => n8587, A2 => n8784, B1 => n7678, B2 => n8582
                           , ZN => n1806);
   U879 : OAI22_X1 port map( A1 => n8587, A2 => n8787, B1 => n7680, B2 => n8582
                           , ZN => n1807);
   U880 : OAI22_X1 port map( A1 => n8628, A2 => n8717, B1 => n7889, B2 => n8627
                           , ZN => n1944);
   U881 : OAI22_X1 port map( A1 => n8628, A2 => n8720, B1 => n7890, B2 => n8627
                           , ZN => n1945);
   U882 : OAI22_X1 port map( A1 => n8628, A2 => n8723, B1 => n7891, B2 => n8627
                           , ZN => n1946);
   U883 : OAI22_X1 port map( A1 => n8628, A2 => n8726, B1 => n7892, B2 => n8627
                           , ZN => n1947);
   U884 : OAI22_X1 port map( A1 => n8628, A2 => n8729, B1 => n7893, B2 => n8627
                           , ZN => n1948);
   U885 : OAI22_X1 port map( A1 => n8629, A2 => n8732, B1 => n7894, B2 => n8627
                           , ZN => n1949);
   U886 : OAI22_X1 port map( A1 => n8629, A2 => n8735, B1 => n7895, B2 => n8627
                           , ZN => n1950);
   U887 : OAI22_X1 port map( A1 => n8629, A2 => n8738, B1 => n7896, B2 => n8627
                           , ZN => n1951);
   U888 : OAI22_X1 port map( A1 => n8629, A2 => n8741, B1 => n7897, B2 => n8627
                           , ZN => n1952);
   U889 : OAI22_X1 port map( A1 => n8629, A2 => n8744, B1 => n7898, B2 => n8627
                           , ZN => n1953);
   U890 : OAI22_X1 port map( A1 => n8630, A2 => n8747, B1 => n7899, B2 => n8627
                           , ZN => n1954);
   U891 : OAI22_X1 port map( A1 => n8630, A2 => n8750, B1 => n7900, B2 => n8627
                           , ZN => n1955);
   U892 : OAI22_X1 port map( A1 => n8630, A2 => n8753, B1 => n7769, B2 => n3167
                           , ZN => n1956);
   U893 : OAI22_X1 port map( A1 => n8630, A2 => n8756, B1 => n7770, B2 => n3167
                           , ZN => n1957);
   U894 : OAI22_X1 port map( A1 => n8630, A2 => n8759, B1 => n7771, B2 => n3167
                           , ZN => n1958);
   U895 : OAI22_X1 port map( A1 => n8631, A2 => n8762, B1 => n7772, B2 => n8627
                           , ZN => n1959);
   U896 : OAI22_X1 port map( A1 => n8631, A2 => n8765, B1 => n7773, B2 => n8627
                           , ZN => n1960);
   U897 : OAI22_X1 port map( A1 => n8631, A2 => n8768, B1 => n7774, B2 => n8627
                           , ZN => n1961);
   U898 : OAI22_X1 port map( A1 => n8631, A2 => n8771, B1 => n7775, B2 => n8627
                           , ZN => n1962);
   U899 : OAI22_X1 port map( A1 => n8631, A2 => n8774, B1 => n7776, B2 => n8627
                           , ZN => n1963);
   U900 : OAI22_X1 port map( A1 => n8632, A2 => n8777, B1 => n7777, B2 => n8627
                           , ZN => n1964);
   U901 : OAI22_X1 port map( A1 => n8632, A2 => n8780, B1 => n7778, B2 => n8627
                           , ZN => n1965);
   U902 : OAI22_X1 port map( A1 => n8632, A2 => n8783, B1 => n7779, B2 => n8627
                           , ZN => n1966);
   U903 : OAI22_X1 port map( A1 => n8632, A2 => n8786, B1 => n7780, B2 => n8627
                           , ZN => n1967);
   U904 : OAI22_X1 port map( A1 => n8646, A2 => n8717, B1 => n7841, B2 => n8645
                           , ZN => n2008);
   U905 : OAI22_X1 port map( A1 => n8646, A2 => n8720, B1 => n7842, B2 => n8645
                           , ZN => n2009);
   U906 : OAI22_X1 port map( A1 => n8646, A2 => n8723, B1 => n7843, B2 => n8645
                           , ZN => n2010);
   U907 : OAI22_X1 port map( A1 => n8646, A2 => n8726, B1 => n7844, B2 => n8645
                           , ZN => n2011);
   U908 : OAI22_X1 port map( A1 => n8646, A2 => n8729, B1 => n7845, B2 => n8645
                           , ZN => n2012);
   U909 : OAI22_X1 port map( A1 => n8647, A2 => n8732, B1 => n7846, B2 => n8645
                           , ZN => n2013);
   U910 : OAI22_X1 port map( A1 => n8647, A2 => n8735, B1 => n7847, B2 => n8645
                           , ZN => n2014);
   U911 : OAI22_X1 port map( A1 => n8647, A2 => n8738, B1 => n7848, B2 => n8645
                           , ZN => n2015);
   U912 : OAI22_X1 port map( A1 => n8647, A2 => n8741, B1 => n7849, B2 => n8645
                           , ZN => n2016);
   U913 : OAI22_X1 port map( A1 => n8647, A2 => n8744, B1 => n7850, B2 => n8645
                           , ZN => n2017);
   U914 : OAI22_X1 port map( A1 => n8648, A2 => n8747, B1 => n7851, B2 => n8645
                           , ZN => n2018);
   U915 : OAI22_X1 port map( A1 => n8648, A2 => n8750, B1 => n7852, B2 => n8645
                           , ZN => n2019);
   U916 : OAI22_X1 port map( A1 => n8648, A2 => n8753, B1 => n7717, B2 => n3164
                           , ZN => n2020);
   U917 : OAI22_X1 port map( A1 => n8648, A2 => n8756, B1 => n7718, B2 => n3164
                           , ZN => n2021);
   U918 : OAI22_X1 port map( A1 => n8648, A2 => n8759, B1 => n7719, B2 => n3164
                           , ZN => n2022);
   U919 : OAI22_X1 port map( A1 => n8649, A2 => n8762, B1 => n7720, B2 => n8645
                           , ZN => n2023);
   U920 : OAI22_X1 port map( A1 => n8649, A2 => n8765, B1 => n7721, B2 => n8645
                           , ZN => n2024);
   U921 : OAI22_X1 port map( A1 => n8649, A2 => n8768, B1 => n7722, B2 => n8645
                           , ZN => n2025);
   U922 : OAI22_X1 port map( A1 => n8649, A2 => n8771, B1 => n7723, B2 => n8645
                           , ZN => n2026);
   U923 : OAI22_X1 port map( A1 => n8649, A2 => n8774, B1 => n7724, B2 => n8645
                           , ZN => n2027);
   U924 : OAI22_X1 port map( A1 => n8650, A2 => n8777, B1 => n7725, B2 => n8645
                           , ZN => n2028);
   U925 : OAI22_X1 port map( A1 => n8650, A2 => n8780, B1 => n7726, B2 => n8645
                           , ZN => n2029);
   U926 : OAI22_X1 port map( A1 => n8650, A2 => n8783, B1 => n7727, B2 => n8645
                           , ZN => n2030);
   U927 : OAI22_X1 port map( A1 => n8650, A2 => n8786, B1 => n7728, B2 => n8645
                           , ZN => n2031);
   U928 : OAI22_X1 port map( A1 => n8655, A2 => n8717, B1 => n7789, B2 => n8654
                           , ZN => n2040);
   U929 : OAI22_X1 port map( A1 => n8655, A2 => n8720, B1 => n7790, B2 => n8654
                           , ZN => n2041);
   U930 : OAI22_X1 port map( A1 => n8655, A2 => n8723, B1 => n7791, B2 => n8654
                           , ZN => n2042);
   U931 : OAI22_X1 port map( A1 => n8655, A2 => n8726, B1 => n7792, B2 => n8654
                           , ZN => n2043);
   U932 : OAI22_X1 port map( A1 => n8655, A2 => n8729, B1 => n7793, B2 => n8654
                           , ZN => n2044);
   U933 : OAI22_X1 port map( A1 => n8656, A2 => n8732, B1 => n7794, B2 => n8654
                           , ZN => n2045);
   U934 : OAI22_X1 port map( A1 => n8656, A2 => n8735, B1 => n7795, B2 => n8654
                           , ZN => n2046);
   U935 : OAI22_X1 port map( A1 => n8656, A2 => n8738, B1 => n7796, B2 => n8654
                           , ZN => n2047);
   U936 : OAI22_X1 port map( A1 => n8656, A2 => n8741, B1 => n7797, B2 => n8654
                           , ZN => n2048);
   U937 : OAI22_X1 port map( A1 => n8656, A2 => n8744, B1 => n7799, B2 => n8654
                           , ZN => n2049);
   U938 : OAI22_X1 port map( A1 => n8657, A2 => n8747, B1 => n7801, B2 => n8654
                           , ZN => n2050);
   U939 : OAI22_X1 port map( A1 => n8657, A2 => n8750, B1 => n7803, B2 => n8654
                           , ZN => n2051);
   U940 : OAI22_X1 port map( A1 => n8657, A2 => n8753, B1 => n7657, B2 => n3162
                           , ZN => n2052);
   U941 : OAI22_X1 port map( A1 => n8657, A2 => n8756, B1 => n7659, B2 => n3162
                           , ZN => n2053);
   U942 : OAI22_X1 port map( A1 => n8657, A2 => n8759, B1 => n7661, B2 => n3162
                           , ZN => n2054);
   U943 : OAI22_X1 port map( A1 => n8658, A2 => n8762, B1 => n7663, B2 => n8654
                           , ZN => n2055);
   U944 : OAI22_X1 port map( A1 => n8658, A2 => n8765, B1 => n7665, B2 => n8654
                           , ZN => n2056);
   U945 : OAI22_X1 port map( A1 => n8658, A2 => n8768, B1 => n7667, B2 => n8654
                           , ZN => n2057);
   U946 : OAI22_X1 port map( A1 => n8658, A2 => n8771, B1 => n7669, B2 => n8654
                           , ZN => n2058);
   U947 : OAI22_X1 port map( A1 => n8658, A2 => n8774, B1 => n7671, B2 => n8654
                           , ZN => n2059);
   U948 : OAI22_X1 port map( A1 => n8659, A2 => n8777, B1 => n7673, B2 => n8654
                           , ZN => n2060);
   U949 : OAI22_X1 port map( A1 => n8659, A2 => n8780, B1 => n7675, B2 => n8654
                           , ZN => n2061);
   U950 : OAI22_X1 port map( A1 => n8659, A2 => n8783, B1 => n7677, B2 => n8654
                           , ZN => n2062);
   U951 : OAI22_X1 port map( A1 => n8659, A2 => n8786, B1 => n7679, B2 => n8654
                           , ZN => n2063);
   U952 : OAI22_X1 port map( A1 => n8664, A2 => n8717, B1 => n8133, B2 => n8663
                           , ZN => n2072);
   U953 : OAI22_X1 port map( A1 => n8664, A2 => n8720, B1 => n8134, B2 => n8663
                           , ZN => n2073);
   U954 : OAI22_X1 port map( A1 => n8664, A2 => n8723, B1 => n8135, B2 => n8663
                           , ZN => n2074);
   U955 : OAI22_X1 port map( A1 => n8664, A2 => n8726, B1 => n8136, B2 => n8663
                           , ZN => n2075);
   U956 : OAI22_X1 port map( A1 => n8664, A2 => n8729, B1 => n8137, B2 => n8663
                           , ZN => n2076);
   U957 : OAI22_X1 port map( A1 => n8665, A2 => n8732, B1 => n8138, B2 => n8663
                           , ZN => n2077);
   U958 : OAI22_X1 port map( A1 => n8665, A2 => n8735, B1 => n8139, B2 => n8663
                           , ZN => n2078);
   U959 : OAI22_X1 port map( A1 => n8665, A2 => n8738, B1 => n8140, B2 => n8663
                           , ZN => n2079);
   U960 : OAI22_X1 port map( A1 => n8665, A2 => n8741, B1 => n8141, B2 => n8663
                           , ZN => n2080);
   U961 : OAI22_X1 port map( A1 => n8665, A2 => n8744, B1 => n8142, B2 => n8663
                           , ZN => n2081);
   U962 : OAI22_X1 port map( A1 => n8666, A2 => n8747, B1 => n8143, B2 => n8663
                           , ZN => n2082);
   U963 : OAI22_X1 port map( A1 => n8666, A2 => n8750, B1 => n8144, B2 => n8663
                           , ZN => n2083);
   U964 : OAI22_X1 port map( A1 => n8666, A2 => n8753, B1 => n8145, B2 => n3160
                           , ZN => n2084);
   U965 : OAI22_X1 port map( A1 => n8666, A2 => n8756, B1 => n8146, B2 => n3160
                           , ZN => n2085);
   U966 : OAI22_X1 port map( A1 => n8666, A2 => n8759, B1 => n8147, B2 => n3160
                           , ZN => n2086);
   U967 : OAI22_X1 port map( A1 => n8667, A2 => n8762, B1 => n8148, B2 => n8663
                           , ZN => n2087);
   U968 : OAI22_X1 port map( A1 => n8667, A2 => n8765, B1 => n8149, B2 => n8663
                           , ZN => n2088);
   U969 : OAI22_X1 port map( A1 => n8667, A2 => n8768, B1 => n8150, B2 => n8663
                           , ZN => n2089);
   U970 : OAI22_X1 port map( A1 => n8667, A2 => n8771, B1 => n8151, B2 => n8663
                           , ZN => n2090);
   U971 : OAI22_X1 port map( A1 => n8667, A2 => n8774, B1 => n8152, B2 => n8663
                           , ZN => n2091);
   U972 : OAI22_X1 port map( A1 => n8668, A2 => n8777, B1 => n8153, B2 => n8663
                           , ZN => n2092);
   U973 : OAI22_X1 port map( A1 => n8668, A2 => n8780, B1 => n8154, B2 => n8663
                           , ZN => n2093);
   U974 : OAI22_X1 port map( A1 => n8668, A2 => n8783, B1 => n8155, B2 => n8663
                           , ZN => n2094);
   U975 : OAI22_X1 port map( A1 => n8668, A2 => n8786, B1 => n8156, B2 => n8663
                           , ZN => n2095);
   U976 : OAI22_X1 port map( A1 => n8691, A2 => n8717, B1 => n7877, B2 => n8690
                           , ZN => n2168);
   U977 : OAI22_X1 port map( A1 => n8691, A2 => n8720, B1 => n7878, B2 => n8690
                           , ZN => n2169);
   U978 : OAI22_X1 port map( A1 => n8691, A2 => n8723, B1 => n7879, B2 => n8690
                           , ZN => n2170);
   U979 : OAI22_X1 port map( A1 => n8691, A2 => n8726, B1 => n7880, B2 => n8690
                           , ZN => n2171);
   U980 : OAI22_X1 port map( A1 => n8691, A2 => n8729, B1 => n7881, B2 => n8690
                           , ZN => n2172);
   U981 : OAI22_X1 port map( A1 => n8692, A2 => n8732, B1 => n7882, B2 => n8690
                           , ZN => n2173);
   U982 : OAI22_X1 port map( A1 => n8692, A2 => n8735, B1 => n7883, B2 => n8690
                           , ZN => n2174);
   U983 : OAI22_X1 port map( A1 => n8692, A2 => n8738, B1 => n7884, B2 => n8690
                           , ZN => n2175);
   U984 : OAI22_X1 port map( A1 => n8692, A2 => n8741, B1 => n7885, B2 => n8690
                           , ZN => n2176);
   U985 : OAI22_X1 port map( A1 => n8692, A2 => n8744, B1 => n7886, B2 => n8690
                           , ZN => n2177);
   U986 : OAI22_X1 port map( A1 => n8693, A2 => n8747, B1 => n7887, B2 => n8690
                           , ZN => n2178);
   U987 : OAI22_X1 port map( A1 => n8693, A2 => n8750, B1 => n7888, B2 => n8690
                           , ZN => n2179);
   U988 : OAI22_X1 port map( A1 => n8693, A2 => n8753, B1 => n7741, B2 => n3154
                           , ZN => n2180);
   U989 : OAI22_X1 port map( A1 => n8693, A2 => n8756, B1 => n7742, B2 => n3154
                           , ZN => n2181);
   U990 : OAI22_X1 port map( A1 => n8693, A2 => n8759, B1 => n7743, B2 => n3154
                           , ZN => n2182);
   U991 : OAI22_X1 port map( A1 => n8694, A2 => n8762, B1 => n7744, B2 => n8690
                           , ZN => n2183);
   U992 : OAI22_X1 port map( A1 => n8694, A2 => n8765, B1 => n7745, B2 => n8690
                           , ZN => n2184);
   U993 : OAI22_X1 port map( A1 => n8694, A2 => n8768, B1 => n7746, B2 => n8690
                           , ZN => n2185);
   U994 : OAI22_X1 port map( A1 => n8694, A2 => n8771, B1 => n7747, B2 => n8690
                           , ZN => n2186);
   U995 : OAI22_X1 port map( A1 => n8694, A2 => n8774, B1 => n7748, B2 => n8690
                           , ZN => n2187);
   U996 : OAI22_X1 port map( A1 => n8695, A2 => n8777, B1 => n7749, B2 => n8690
                           , ZN => n2188);
   U997 : OAI22_X1 port map( A1 => n8695, A2 => n8780, B1 => n7750, B2 => n8690
                           , ZN => n2189);
   U998 : OAI22_X1 port map( A1 => n8695, A2 => n8783, B1 => n7751, B2 => n8690
                           , ZN => n2190);
   U999 : OAI22_X1 port map( A1 => n8695, A2 => n8786, B1 => n7752, B2 => n8690
                           , ZN => n2191);
   U1000 : OAI22_X1 port map( A1 => n8700, A2 => n8717, B1 => n7729, B2 => 
                           n8699, ZN => n2200);
   U1001 : OAI22_X1 port map( A1 => n8700, A2 => n8720, B1 => n7730, B2 => 
                           n8699, ZN => n2201);
   U1002 : OAI22_X1 port map( A1 => n8700, A2 => n8723, B1 => n7731, B2 => 
                           n8699, ZN => n2202);
   U1003 : OAI22_X1 port map( A1 => n8700, A2 => n8726, B1 => n7732, B2 => 
                           n8699, ZN => n2203);
   U1004 : OAI22_X1 port map( A1 => n8700, A2 => n8729, B1 => n7733, B2 => 
                           n8699, ZN => n2204);
   U1005 : OAI22_X1 port map( A1 => n8701, A2 => n8732, B1 => n7734, B2 => 
                           n8699, ZN => n2205);
   U1006 : OAI22_X1 port map( A1 => n8701, A2 => n8735, B1 => n7735, B2 => 
                           n8699, ZN => n2206);
   U1007 : OAI22_X1 port map( A1 => n8701, A2 => n8738, B1 => n7736, B2 => 
                           n8699, ZN => n2207);
   U1008 : OAI22_X1 port map( A1 => n8701, A2 => n8741, B1 => n7737, B2 => 
                           n8699, ZN => n2208);
   U1009 : OAI22_X1 port map( A1 => n8701, A2 => n8744, B1 => n7738, B2 => 
                           n8699, ZN => n2209);
   U1010 : OAI22_X1 port map( A1 => n8702, A2 => n8747, B1 => n7739, B2 => 
                           n8699, ZN => n2210);
   U1011 : OAI22_X1 port map( A1 => n8702, A2 => n8750, B1 => n7740, B2 => 
                           n8699, ZN => n2211);
   U1012 : OAI22_X1 port map( A1 => n8702, A2 => n8753, B1 => n7645, B2 => 
                           n3152, ZN => n2212);
   U1013 : OAI22_X1 port map( A1 => n8702, A2 => n8756, B1 => n7646, B2 => 
                           n3152, ZN => n2213);
   U1014 : OAI22_X1 port map( A1 => n8702, A2 => n8759, B1 => n7647, B2 => 
                           n3152, ZN => n2214);
   U1015 : OAI22_X1 port map( A1 => n8703, A2 => n8762, B1 => n7648, B2 => 
                           n8699, ZN => n2215);
   U1016 : OAI22_X1 port map( A1 => n8703, A2 => n8765, B1 => n7649, B2 => 
                           n8699, ZN => n2216);
   U1017 : OAI22_X1 port map( A1 => n8703, A2 => n8768, B1 => n7650, B2 => 
                           n8699, ZN => n2217);
   U1018 : OAI22_X1 port map( A1 => n8703, A2 => n8771, B1 => n7651, B2 => 
                           n8699, ZN => n2218);
   U1019 : OAI22_X1 port map( A1 => n8703, A2 => n8774, B1 => n7652, B2 => 
                           n8699, ZN => n2219);
   U1020 : OAI22_X1 port map( A1 => n8704, A2 => n8777, B1 => n7653, B2 => 
                           n8699, ZN => n2220);
   U1021 : OAI22_X1 port map( A1 => n8704, A2 => n8780, B1 => n7654, B2 => 
                           n8699, ZN => n2221);
   U1022 : OAI22_X1 port map( A1 => n8704, A2 => n8783, B1 => n7655, B2 => 
                           n8699, ZN => n2222);
   U1023 : OAI22_X1 port map( A1 => n8704, A2 => n8786, B1 => n7656, B2 => 
                           n8699, ZN => n2223);
   U1024 : OAI22_X1 port map( A1 => n8709, A2 => n8717, B1 => n8109, B2 => 
                           n8708, ZN => n2232);
   U1025 : OAI22_X1 port map( A1 => n8709, A2 => n8720, B1 => n8110, B2 => 
                           n8708, ZN => n2233);
   U1026 : OAI22_X1 port map( A1 => n8709, A2 => n8723, B1 => n8111, B2 => 
                           n8708, ZN => n2234);
   U1027 : OAI22_X1 port map( A1 => n8709, A2 => n8726, B1 => n8112, B2 => 
                           n8708, ZN => n2235);
   U1028 : OAI22_X1 port map( A1 => n8709, A2 => n8729, B1 => n8113, B2 => 
                           n8708, ZN => n2236);
   U1029 : OAI22_X1 port map( A1 => n8710, A2 => n8732, B1 => n8114, B2 => 
                           n8708, ZN => n2237);
   U1030 : OAI22_X1 port map( A1 => n8710, A2 => n8735, B1 => n8115, B2 => 
                           n8708, ZN => n2238);
   U1031 : OAI22_X1 port map( A1 => n8710, A2 => n8738, B1 => n8116, B2 => 
                           n8708, ZN => n2239);
   U1032 : OAI22_X1 port map( A1 => n8710, A2 => n8741, B1 => n8117, B2 => 
                           n8708, ZN => n2240);
   U1033 : OAI22_X1 port map( A1 => n8710, A2 => n8744, B1 => n8118, B2 => 
                           n8708, ZN => n2241);
   U1034 : OAI22_X1 port map( A1 => n8711, A2 => n8747, B1 => n8119, B2 => 
                           n8708, ZN => n2242);
   U1035 : OAI22_X1 port map( A1 => n8711, A2 => n8750, B1 => n8120, B2 => 
                           n8708, ZN => n2243);
   U1036 : OAI22_X1 port map( A1 => n8711, A2 => n8753, B1 => n8121, B2 => 
                           n3150, ZN => n2244);
   U1037 : OAI22_X1 port map( A1 => n8711, A2 => n8756, B1 => n8122, B2 => 
                           n3150, ZN => n2245);
   U1038 : OAI22_X1 port map( A1 => n8711, A2 => n8759, B1 => n8123, B2 => 
                           n3150, ZN => n2246);
   U1039 : OAI22_X1 port map( A1 => n8712, A2 => n8762, B1 => n8124, B2 => 
                           n8708, ZN => n2247);
   U1040 : OAI22_X1 port map( A1 => n8712, A2 => n8765, B1 => n8125, B2 => 
                           n8708, ZN => n2248);
   U1041 : OAI22_X1 port map( A1 => n8712, A2 => n8768, B1 => n8126, B2 => 
                           n8708, ZN => n2249);
   U1042 : OAI22_X1 port map( A1 => n8712, A2 => n8771, B1 => n8127, B2 => 
                           n8708, ZN => n2250);
   U1043 : OAI22_X1 port map( A1 => n8712, A2 => n8774, B1 => n8128, B2 => 
                           n8708, ZN => n2251);
   U1044 : OAI22_X1 port map( A1 => n8713, A2 => n8777, B1 => n8129, B2 => 
                           n8708, ZN => n2252);
   U1045 : OAI22_X1 port map( A1 => n8713, A2 => n8780, B1 => n8130, B2 => 
                           n8708, ZN => n2253);
   U1046 : OAI22_X1 port map( A1 => n8713, A2 => n8783, B1 => n8131, B2 => 
                           n8708, ZN => n2254);
   U1047 : OAI22_X1 port map( A1 => n8713, A2 => n8786, B1 => n8132, B2 => 
                           n8708, ZN => n2255);
   U1048 : OAI22_X1 port map( A1 => n8811, A2 => n8717, B1 => n8181, B2 => 
                           n8810, ZN => n2264);
   U1049 : OAI22_X1 port map( A1 => n8811, A2 => n8720, B1 => n8182, B2 => 
                           n8810, ZN => n2265);
   U1050 : OAI22_X1 port map( A1 => n8811, A2 => n8723, B1 => n8183, B2 => 
                           n8810, ZN => n2266);
   U1051 : OAI22_X1 port map( A1 => n8811, A2 => n8726, B1 => n8184, B2 => 
                           n8810, ZN => n2267);
   U1052 : OAI22_X1 port map( A1 => n8811, A2 => n8729, B1 => n8185, B2 => 
                           n8810, ZN => n2268);
   U1053 : OAI22_X1 port map( A1 => n8812, A2 => n8732, B1 => n8186, B2 => 
                           n8810, ZN => n2269);
   U1054 : OAI22_X1 port map( A1 => n8812, A2 => n8735, B1 => n8187, B2 => 
                           n8810, ZN => n2270);
   U1055 : OAI22_X1 port map( A1 => n8812, A2 => n8738, B1 => n8188, B2 => 
                           n8810, ZN => n2271);
   U1056 : OAI22_X1 port map( A1 => n8812, A2 => n8741, B1 => n8189, B2 => 
                           n8810, ZN => n2272);
   U1057 : OAI22_X1 port map( A1 => n8812, A2 => n8744, B1 => n8190, B2 => 
                           n8810, ZN => n2273);
   U1058 : OAI22_X1 port map( A1 => n8813, A2 => n8747, B1 => n8191, B2 => 
                           n8810, ZN => n2274);
   U1059 : OAI22_X1 port map( A1 => n8813, A2 => n8750, B1 => n8192, B2 => 
                           n8810, ZN => n2275);
   U1060 : OAI22_X1 port map( A1 => n8813, A2 => n8753, B1 => n8193, B2 => 
                           n3116, ZN => n2276);
   U1061 : OAI22_X1 port map( A1 => n8813, A2 => n8756, B1 => n8194, B2 => 
                           n3116, ZN => n2277);
   U1062 : OAI22_X1 port map( A1 => n8813, A2 => n8759, B1 => n8195, B2 => 
                           n3116, ZN => n2278);
   U1063 : OAI22_X1 port map( A1 => n8814, A2 => n8762, B1 => n8196, B2 => 
                           n8810, ZN => n2279);
   U1064 : OAI22_X1 port map( A1 => n8814, A2 => n8765, B1 => n8197, B2 => 
                           n8810, ZN => n2280);
   U1065 : OAI22_X1 port map( A1 => n8814, A2 => n8768, B1 => n8198, B2 => 
                           n8810, ZN => n2281);
   U1066 : OAI22_X1 port map( A1 => n8814, A2 => n8771, B1 => n8199, B2 => 
                           n8810, ZN => n2282);
   U1067 : OAI22_X1 port map( A1 => n8814, A2 => n8774, B1 => n8200, B2 => 
                           n8810, ZN => n2283);
   U1068 : OAI22_X1 port map( A1 => n8815, A2 => n8777, B1 => n8201, B2 => 
                           n8810, ZN => n2284);
   U1069 : OAI22_X1 port map( A1 => n8815, A2 => n8780, B1 => n8202, B2 => 
                           n8810, ZN => n2285);
   U1070 : OAI22_X1 port map( A1 => n8815, A2 => n8783, B1 => n8203, B2 => 
                           n8810, ZN => n2286);
   U1071 : OAI22_X1 port map( A1 => n8815, A2 => n8786, B1 => n8204, B2 => 
                           n8810, ZN => n2287);
   U1072 : NOR3_X1 port map( A1 => n845, A2 => ADD_RD2(4), A3 => n846, ZN => 
                           n2489);
   U1073 : NOR3_X1 port map( A1 => n844, A2 => n845, A3 => n846, ZN => n2471);
   U1074 : NOR3_X1 port map( A1 => n839, A2 => n840, A3 => n841, ZN => n3103);
   U1075 : NOR3_X1 port map( A1 => n840, A2 => ADD_RD1(4), A3 => n841, ZN => 
                           n3094);
   U1076 : NAND2_X1 port map( A1 => n3095, A2 => n3112, ZN => n2533);
   U1077 : NAND2_X1 port map( A1 => n3096, A2 => n3112, ZN => n2529);
   U1078 : NAND2_X1 port map( A1 => n3096, A2 => n3105, ZN => n2527);
   U1079 : NAND2_X1 port map( A1 => n3099, A2 => n3112, ZN => n2532);
   U1080 : BUF_X1 port map( A => n833, Z => n9024);
   U1081 : BUF_X1 port map( A => n833, Z => n9023);
   U1082 : NAND2_X1 port map( A1 => n2475, A2 => n2474, ZN => n896);
   U1083 : NAND2_X1 port map( A1 => n2475, A2 => n2476, ZN => n855);
   U1084 : BUF_X1 port map( A => n884, Z => n8957);
   U1085 : BUF_X1 port map( A => n2506, Z => n8909);
   U1086 : BUF_X1 port map( A => n833, Z => n9021);
   U1087 : BUF_X1 port map( A => n833, Z => n9020);
   U1088 : BUF_X1 port map( A => n3147, Z => n8718);
   U1089 : BUF_X1 port map( A => n3146, Z => n8721);
   U1090 : BUF_X1 port map( A => n3145, Z => n8724);
   U1091 : BUF_X1 port map( A => n3144, Z => n8727);
   U1092 : BUF_X1 port map( A => n3143, Z => n8730);
   U1093 : BUF_X1 port map( A => n3142, Z => n8733);
   U1094 : BUF_X1 port map( A => n3141, Z => n8736);
   U1095 : BUF_X1 port map( A => n3140, Z => n8739);
   U1096 : BUF_X1 port map( A => n3139, Z => n8742);
   U1097 : BUF_X1 port map( A => n3138, Z => n8745);
   U1098 : BUF_X1 port map( A => n3137, Z => n8748);
   U1099 : BUF_X1 port map( A => n3136, Z => n8751);
   U1100 : BUF_X1 port map( A => n3135, Z => n8754);
   U1101 : BUF_X1 port map( A => n3134, Z => n8757);
   U1102 : BUF_X1 port map( A => n3133, Z => n8760);
   U1103 : BUF_X1 port map( A => n3132, Z => n8763);
   U1104 : BUF_X1 port map( A => n3131, Z => n8766);
   U1105 : BUF_X1 port map( A => n3130, Z => n8769);
   U1106 : BUF_X1 port map( A => n3129, Z => n8772);
   U1107 : BUF_X1 port map( A => n3128, Z => n8775);
   U1108 : BUF_X1 port map( A => n3127, Z => n8778);
   U1109 : BUF_X1 port map( A => n3126, Z => n8781);
   U1110 : BUF_X1 port map( A => n3125, Z => n8784);
   U1111 : BUF_X1 port map( A => n3124, Z => n8787);
   U1112 : BUF_X1 port map( A => n3123, Z => n8790);
   U1113 : BUF_X1 port map( A => n3122, Z => n8793);
   U1114 : BUF_X1 port map( A => n3121, Z => n8796);
   U1115 : BUF_X1 port map( A => n3120, Z => n8799);
   U1116 : BUF_X1 port map( A => n3119, Z => n8802);
   U1117 : BUF_X1 port map( A => n3118, Z => n8805);
   U1118 : BUF_X1 port map( A => n3117, Z => n8808);
   U1119 : BUF_X1 port map( A => n3115, Z => n8820);
   U1120 : BUF_X1 port map( A => n3147, Z => n8717);
   U1121 : BUF_X1 port map( A => n3146, Z => n8720);
   U1122 : BUF_X1 port map( A => n3145, Z => n8723);
   U1123 : BUF_X1 port map( A => n3144, Z => n8726);
   U1124 : BUF_X1 port map( A => n3143, Z => n8729);
   U1125 : BUF_X1 port map( A => n3142, Z => n8732);
   U1126 : BUF_X1 port map( A => n3141, Z => n8735);
   U1127 : BUF_X1 port map( A => n3140, Z => n8738);
   U1128 : BUF_X1 port map( A => n3139, Z => n8741);
   U1129 : BUF_X1 port map( A => n3138, Z => n8744);
   U1130 : BUF_X1 port map( A => n3137, Z => n8747);
   U1131 : BUF_X1 port map( A => n3136, Z => n8750);
   U1132 : BUF_X1 port map( A => n3135, Z => n8753);
   U1133 : BUF_X1 port map( A => n3134, Z => n8756);
   U1134 : BUF_X1 port map( A => n3133, Z => n8759);
   U1135 : BUF_X1 port map( A => n3132, Z => n8762);
   U1136 : BUF_X1 port map( A => n3131, Z => n8765);
   U1137 : BUF_X1 port map( A => n3130, Z => n8768);
   U1138 : BUF_X1 port map( A => n3129, Z => n8771);
   U1139 : BUF_X1 port map( A => n3128, Z => n8774);
   U1140 : BUF_X1 port map( A => n3127, Z => n8777);
   U1141 : BUF_X1 port map( A => n3126, Z => n8780);
   U1142 : BUF_X1 port map( A => n3125, Z => n8783);
   U1143 : BUF_X1 port map( A => n3124, Z => n8786);
   U1144 : BUF_X1 port map( A => n3123, Z => n8789);
   U1145 : BUF_X1 port map( A => n3122, Z => n8792);
   U1146 : BUF_X1 port map( A => n3121, Z => n8795);
   U1147 : BUF_X1 port map( A => n3120, Z => n8798);
   U1148 : BUF_X1 port map( A => n3119, Z => n8801);
   U1149 : BUF_X1 port map( A => n3118, Z => n8804);
   U1150 : BUF_X1 port map( A => n3117, Z => n8807);
   U1151 : BUF_X1 port map( A => n3115, Z => n8819);
   U1152 : NAND2_X1 port map( A1 => n2473, A2 => n2474, ZN => n856);
   U1153 : NAND2_X1 port map( A1 => n2473, A2 => n2482, ZN => n865);
   U1154 : BUF_X1 port map( A => n833, Z => n9022);
   U1155 : NAND2_X1 port map( A1 => n3102, A2 => n3107, ZN => n2518);
   U1156 : BUF_X1 port map( A => n884, Z => n8958);
   U1157 : BUF_X1 port map( A => n2506, Z => n8910);
   U1158 : BUF_X1 port map( A => n3147, Z => n8719);
   U1159 : BUF_X1 port map( A => n3146, Z => n8722);
   U1160 : BUF_X1 port map( A => n3145, Z => n8725);
   U1161 : BUF_X1 port map( A => n3144, Z => n8728);
   U1162 : BUF_X1 port map( A => n3143, Z => n8731);
   U1163 : BUF_X1 port map( A => n3142, Z => n8734);
   U1164 : BUF_X1 port map( A => n3141, Z => n8737);
   U1165 : BUF_X1 port map( A => n3140, Z => n8740);
   U1166 : BUF_X1 port map( A => n3139, Z => n8743);
   U1167 : BUF_X1 port map( A => n3138, Z => n8746);
   U1168 : BUF_X1 port map( A => n3137, Z => n8749);
   U1169 : BUF_X1 port map( A => n3136, Z => n8752);
   U1170 : BUF_X1 port map( A => n3135, Z => n8755);
   U1171 : BUF_X1 port map( A => n3134, Z => n8758);
   U1172 : BUF_X1 port map( A => n3133, Z => n8761);
   U1173 : BUF_X1 port map( A => n3132, Z => n8764);
   U1174 : BUF_X1 port map( A => n3131, Z => n8767);
   U1175 : BUF_X1 port map( A => n3130, Z => n8770);
   U1176 : BUF_X1 port map( A => n3129, Z => n8773);
   U1177 : BUF_X1 port map( A => n3128, Z => n8776);
   U1178 : BUF_X1 port map( A => n3127, Z => n8779);
   U1179 : BUF_X1 port map( A => n3126, Z => n8782);
   U1180 : BUF_X1 port map( A => n3125, Z => n8785);
   U1181 : BUF_X1 port map( A => n3124, Z => n8788);
   U1182 : BUF_X1 port map( A => n3123, Z => n8791);
   U1183 : BUF_X1 port map( A => n3122, Z => n8794);
   U1184 : BUF_X1 port map( A => n3121, Z => n8797);
   U1185 : BUF_X1 port map( A => n3120, Z => n8800);
   U1186 : BUF_X1 port map( A => n3119, Z => n8803);
   U1187 : BUF_X1 port map( A => n3118, Z => n8806);
   U1188 : BUF_X1 port map( A => n3117, Z => n8809);
   U1189 : BUF_X1 port map( A => n3115, Z => n8821);
   U1190 : NAND2_X1 port map( A1 => n3097, A2 => n3095, ZN => n2502);
   U1191 : NAND2_X1 port map( A1 => n3105, A2 => n3095, ZN => n2534);
   U1192 : NAND2_X1 port map( A1 => n3106, A2 => n3095, ZN => n2526);
   U1193 : NAND2_X1 port map( A1 => n3107, A2 => n3095, ZN => n2530);
   U1194 : NAND2_X1 port map( A1 => n3103, A2 => n3095, ZN => n2544);
   U1195 : NAND2_X1 port map( A1 => n3100, A2 => n3096, ZN => n2507);
   U1196 : NAND2_X1 port map( A1 => n3094, A2 => n3096, ZN => n2503);
   U1197 : NAND2_X1 port map( A1 => n3106, A2 => n3096, ZN => n2539);
   U1198 : NAND2_X1 port map( A1 => n3097, A2 => n3096, ZN => n2543);
   U1199 : NAND2_X1 port map( A1 => n2491, A2 => n2480, ZN => n885);
   U1200 : NAND2_X1 port map( A1 => n2479, A2 => n2480, ZN => n880);
   U1201 : NAND2_X1 port map( A1 => n2474, A2 => n2480, ZN => n871);
   U1202 : NAND2_X1 port map( A1 => n2471, A2 => n2480, ZN => n860);
   U1203 : NAND2_X1 port map( A1 => n2478, A2 => n2480, ZN => n866);
   U1204 : NAND2_X1 port map( A1 => n3097, A2 => n3099, ZN => n2508);
   U1205 : NAND2_X1 port map( A1 => n3105, A2 => n3099, ZN => n2528);
   U1206 : NAND2_X1 port map( A1 => n3107, A2 => n3099, ZN => n2531);
   U1207 : NAND2_X1 port map( A1 => n3106, A2 => n3099, ZN => n2538);
   U1208 : NAND2_X1 port map( A1 => n2491, A2 => n2475, ZN => n890);
   U1209 : NAND2_X1 port map( A1 => n2474, A2 => n2472, ZN => n870);
   U1210 : NAND2_X1 port map( A1 => n2489, A2 => n2473, ZN => n881);
   U1211 : NAND2_X1 port map( A1 => n2479, A2 => n2473, ZN => n861);
   U1212 : NAND2_X1 port map( A1 => n3100, A2 => n3102, ZN => n2512);
   U1213 : BUF_X1 port map( A => n884, Z => n8959);
   U1214 : BUF_X1 port map( A => n2506, Z => n8911);
   U1215 : NAND2_X1 port map( A1 => n2489, A2 => n2472, ZN => n886);
   U1216 : INV_X1 port map( A => ADD_RD2(4), ZN => n844);
   U1217 : INV_X1 port map( A => ADD_RD1(4), ZN => n839);
   U1218 : AND2_X1 port map( A1 => n3096, A2 => n3107, ZN => n2541);
   U1219 : AND2_X1 port map( A1 => n2480, A2 => n2476, ZN => n874);
   U1220 : AND2_X1 port map( A1 => n2475, A2 => n2479, ZN => n893);
   U1221 : AND2_X1 port map( A1 => n2475, A2 => n2478, ZN => n898);
   U1222 : AND2_X1 port map( A1 => n2475, A2 => n2482, ZN => n899);
   U1223 : AND2_X1 port map( A1 => n2473, A2 => n2476, ZN => n868);
   U1224 : AND2_X1 port map( A1 => n3102, A2 => n3097, ZN => n2515);
   U1225 : AND2_X1 port map( A1 => n3102, A2 => n3106, ZN => n2520);
   U1226 : AND2_X1 port map( A1 => n3102, A2 => n3105, ZN => n2521);
   U1227 : AND2_X1 port map( A1 => n3102, A2 => n3112, ZN => n2540);
   U1228 : AND2_X1 port map( A1 => n2472, A2 => n2476, ZN => n875);
   U1229 : AND2_X1 port map( A1 => n3100, A2 => n3095, ZN => n2510);
   U1230 : AND2_X1 port map( A1 => n3094, A2 => n3095, ZN => n2505);
   U1231 : AND2_X1 port map( A1 => n3103, A2 => n3096, ZN => n2535);
   U1232 : AND2_X1 port map( A1 => n2489, A2 => n2480, ZN => n883);
   U1233 : AND2_X1 port map( A1 => n2482, A2 => n2480, ZN => n873);
   U1234 : AND2_X1 port map( A1 => n3094, A2 => n3099, ZN => n2511);
   U1235 : AND2_X1 port map( A1 => n3100, A2 => n3099, ZN => n2516);
   U1236 : AND2_X1 port map( A1 => n3103, A2 => n3099, ZN => n2536);
   U1237 : AND2_X1 port map( A1 => n2491, A2 => n2473, ZN => n888);
   U1238 : AND2_X1 port map( A1 => n2471, A2 => n2473, ZN => n858);
   U1239 : AND2_X1 port map( A1 => n2478, A2 => n2473, ZN => n863);
   U1240 : AND2_X1 port map( A1 => n2479, A2 => n2472, ZN => n889);
   U1241 : AND2_X1 port map( A1 => n2491, A2 => n2472, ZN => n894);
   U1242 : AND2_X1 port map( A1 => n2471, A2 => n2472, ZN => n859);
   U1243 : AND2_X1 port map( A1 => n2478, A2 => n2472, ZN => n864);
   U1244 : AND2_X1 port map( A1 => n2482, A2 => n2472, ZN => n869);
   U1245 : BUF_X1 port map( A => n3190, Z => n8437);
   U1246 : OAI21_X1 port map( B1 => n3163, B2 => n3183, A => n9024, ZN => n3190
                           );
   U1247 : INV_X1 port map( A => ADD_WR(4), ZN => n834);
   U1248 : INV_X1 port map( A => n3162, ZN => n8662);
   U1249 : OAI21_X1 port map( B1 => n3148, B2 => n3163, A => n9024, ZN => n3162
                           );
   U1250 : INV_X1 port map( A => n3160, ZN => n8671);
   U1251 : OAI21_X1 port map( B1 => n3148, B2 => n3161, A => n9024, ZN => n3160
                           );
   U1252 : INV_X1 port map( A => n3158, ZN => n8680);
   U1253 : OAI21_X1 port map( B1 => n3148, B2 => n3159, A => n9024, ZN => n3158
                           );
   U1254 : INV_X1 port map( A => n3156, ZN => n8689);
   U1255 : OAI21_X1 port map( B1 => n3148, B2 => n3157, A => n9024, ZN => n3156
                           );
   U1256 : INV_X1 port map( A => n3154, ZN => n8698);
   U1257 : OAI21_X1 port map( B1 => n3148, B2 => n3155, A => n9024, ZN => n3154
                           );
   U1258 : INV_X1 port map( A => n3152, ZN => n8707);
   U1259 : OAI21_X1 port map( B1 => n3148, B2 => n3153, A => n9024, ZN => n3152
                           );
   U1260 : INV_X1 port map( A => n3150, ZN => n8716);
   U1261 : OAI21_X1 port map( B1 => n3148, B2 => n3151, A => n9025, ZN => n3150
                           );
   U1262 : INV_X1 port map( A => n3116, ZN => n8818);
   U1263 : OAI21_X1 port map( B1 => n3148, B2 => n3149, A => n9025, ZN => n3116
                           );
   U1264 : INV_X1 port map( A => n3189, ZN => n8455);
   U1265 : OAI21_X1 port map( B1 => n3161, B2 => n3183, A => n9022, ZN => n3189
                           );
   U1266 : INV_X1 port map( A => n3188, ZN => n8464);
   U1267 : OAI21_X1 port map( B1 => n3159, B2 => n3183, A => n9022, ZN => n3188
                           );
   U1268 : INV_X1 port map( A => n3187, ZN => n8473);
   U1269 : OAI21_X1 port map( B1 => n3157, B2 => n3183, A => n9022, ZN => n3187
                           );
   U1270 : INV_X1 port map( A => n3186, ZN => n8482);
   U1271 : OAI21_X1 port map( B1 => n3155, B2 => n3183, A => n9023, ZN => n3186
                           );
   U1272 : INV_X1 port map( A => n3185, ZN => n8491);
   U1273 : OAI21_X1 port map( B1 => n3153, B2 => n3183, A => n9022, ZN => n3185
                           );
   U1274 : INV_X1 port map( A => n3184, ZN => n8500);
   U1275 : OAI21_X1 port map( B1 => n3151, B2 => n3183, A => n9023, ZN => n3184
                           );
   U1276 : INV_X1 port map( A => n3182, ZN => n8509);
   U1277 : OAI21_X1 port map( B1 => n3149, B2 => n3183, A => n9023, ZN => n3182
                           );
   U1278 : INV_X1 port map( A => n3181, ZN => n8518);
   U1279 : OAI21_X1 port map( B1 => n3163, B2 => n3174, A => n9023, ZN => n3181
                           );
   U1280 : INV_X1 port map( A => n3180, ZN => n8527);
   U1281 : OAI21_X1 port map( B1 => n3161, B2 => n3174, A => n9023, ZN => n3180
                           );
   U1282 : INV_X1 port map( A => n3179, ZN => n8536);
   U1283 : OAI21_X1 port map( B1 => n3159, B2 => n3174, A => n9023, ZN => n3179
                           );
   U1284 : INV_X1 port map( A => n3178, ZN => n8545);
   U1285 : OAI21_X1 port map( B1 => n3157, B2 => n3174, A => n9023, ZN => n3178
                           );
   U1286 : INV_X1 port map( A => n3177, ZN => n8554);
   U1287 : OAI21_X1 port map( B1 => n3155, B2 => n3174, A => n9023, ZN => n3177
                           );
   U1288 : INV_X1 port map( A => n3176, ZN => n8563);
   U1289 : OAI21_X1 port map( B1 => n3153, B2 => n3174, A => n9023, ZN => n3176
                           );
   U1290 : INV_X1 port map( A => n3175, ZN => n8572);
   U1291 : OAI21_X1 port map( B1 => n3151, B2 => n3174, A => n9023, ZN => n3175
                           );
   U1292 : INV_X1 port map( A => n3173, ZN => n8581);
   U1293 : OAI21_X1 port map( B1 => n3149, B2 => n3174, A => n9023, ZN => n3173
                           );
   U1294 : INV_X1 port map( A => n3172, ZN => n8590);
   U1295 : OAI21_X1 port map( B1 => n3163, B2 => n3165, A => n9023, ZN => n3172
                           );
   U1296 : INV_X1 port map( A => n3171, ZN => n8599);
   U1297 : OAI21_X1 port map( B1 => n3161, B2 => n3165, A => n9023, ZN => n3171
                           );
   U1298 : INV_X1 port map( A => n3170, ZN => n8608);
   U1299 : OAI21_X1 port map( B1 => n3159, B2 => n3165, A => n9024, ZN => n3170
                           );
   U1300 : INV_X1 port map( A => n3169, ZN => n8617);
   U1301 : OAI21_X1 port map( B1 => n3157, B2 => n3165, A => n9024, ZN => n3169
                           );
   U1302 : INV_X1 port map( A => n3168, ZN => n8626);
   U1303 : OAI21_X1 port map( B1 => n3155, B2 => n3165, A => n9024, ZN => n3168
                           );
   U1304 : INV_X1 port map( A => n3167, ZN => n8635);
   U1305 : OAI21_X1 port map( B1 => n3153, B2 => n3165, A => n9024, ZN => n3167
                           );
   U1306 : INV_X1 port map( A => n3166, ZN => n8644);
   U1307 : OAI21_X1 port map( B1 => n3151, B2 => n3165, A => n9024, ZN => n3166
                           );
   U1308 : INV_X1 port map( A => n3164, ZN => n8653);
   U1309 : OAI21_X1 port map( B1 => n3149, B2 => n3165, A => n9024, ZN => n3164
                           );
   U1310 : OAI221_X1 port map( B1 => n6883, B2 => n8982, C1 => n6691, C2 => 
                           n8979, A => n1035, ZN => n1028);
   U1311 : AOI222_X1 port map( A1 => n3655, A2 => n8976, B1 => n6579, B2 => 
                           n8973, C1 => n3847, C2 => n8970, ZN => n1035);
   U1312 : OAI221_X1 port map( B1 => n6884, B2 => n8982, C1 => n6692, C2 => 
                           n8979, A => n1053, ZN => n1046);
   U1313 : AOI222_X1 port map( A1 => n3656, A2 => n8976, B1 => n6580, B2 => 
                           n8973, C1 => n3848, C2 => n8970, ZN => n1053);
   U1314 : OAI221_X1 port map( B1 => n6885, B2 => n8982, C1 => n6693, C2 => 
                           n8979, A => n1071, ZN => n1064);
   U1315 : AOI222_X1 port map( A1 => n3657, A2 => n8976, B1 => n6581, B2 => 
                           n8973, C1 => n3849, C2 => n8970, ZN => n1071);
   U1316 : OAI221_X1 port map( B1 => n6886, B2 => n8982, C1 => n6694, C2 => 
                           n8979, A => n1089, ZN => n1082);
   U1317 : AOI222_X1 port map( A1 => n3658, A2 => n8976, B1 => n6582, B2 => 
                           n8973, C1 => n3850, C2 => n8970, ZN => n1089);
   U1318 : OAI221_X1 port map( B1 => n6887, B2 => n8982, C1 => n6695, C2 => 
                           n8979, A => n1107, ZN => n1100);
   U1319 : AOI222_X1 port map( A1 => n3659, A2 => n8976, B1 => n6583, B2 => 
                           n8973, C1 => n3851, C2 => n8970, ZN => n1107);
   U1320 : OAI221_X1 port map( B1 => n6888, B2 => n8982, C1 => n6696, C2 => 
                           n8979, A => n1125, ZN => n1118);
   U1321 : AOI222_X1 port map( A1 => n3660, A2 => n8976, B1 => n6584, B2 => 
                           n8973, C1 => n3852, C2 => n8970, ZN => n1125);
   U1322 : OAI221_X1 port map( B1 => n6889, B2 => n8982, C1 => n6697, C2 => 
                           n8979, A => n1143, ZN => n1136);
   U1323 : AOI222_X1 port map( A1 => n3661, A2 => n8976, B1 => n6585, B2 => 
                           n8973, C1 => n3853, C2 => n8970, ZN => n1143);
   U1324 : OAI221_X1 port map( B1 => n6890, B2 => n8982, C1 => n6698, C2 => 
                           n8979, A => n1161, ZN => n1154);
   U1325 : AOI222_X1 port map( A1 => n3662, A2 => n8976, B1 => n6586, B2 => 
                           n8973, C1 => n3854, C2 => n8970, ZN => n1161);
   U1326 : OAI221_X1 port map( B1 => n6891, B2 => n8982, C1 => n6699, C2 => 
                           n8979, A => n1179, ZN => n1172);
   U1327 : AOI222_X1 port map( A1 => n3663, A2 => n8976, B1 => n6587, B2 => 
                           n8973, C1 => n3855, C2 => n8970, ZN => n1179);
   U1328 : OAI221_X1 port map( B1 => n6892, B2 => n8982, C1 => n6700, C2 => 
                           n8979, A => n1197, ZN => n1190);
   U1329 : AOI222_X1 port map( A1 => n3664, A2 => n8976, B1 => n6588, B2 => 
                           n8973, C1 => n3856, C2 => n8970, ZN => n1197);
   U1330 : OAI221_X1 port map( B1 => n6893, B2 => n8982, C1 => n6701, C2 => 
                           n8979, A => n1215, ZN => n1208);
   U1331 : AOI222_X1 port map( A1 => n3665, A2 => n8976, B1 => n6589, B2 => 
                           n8973, C1 => n3857, C2 => n8970, ZN => n1215);
   U1332 : OAI221_X1 port map( B1 => n6894, B2 => n8982, C1 => n6702, C2 => 
                           n8979, A => n1233, ZN => n1226);
   U1333 : AOI222_X1 port map( A1 => n3666, A2 => n8976, B1 => n6590, B2 => 
                           n8973, C1 => n3858, C2 => n8970, ZN => n1233);
   U1334 : OAI221_X1 port map( B1 => n6895, B2 => n8981, C1 => n6703, C2 => 
                           n8978, A => n1251, ZN => n1244);
   U1335 : AOI222_X1 port map( A1 => n3667, A2 => n8975, B1 => n6591, B2 => 
                           n8972, C1 => n3859, C2 => n8969, ZN => n1251);
   U1336 : OAI221_X1 port map( B1 => n6896, B2 => n8981, C1 => n6704, C2 => 
                           n8978, A => n1269, ZN => n1262);
   U1337 : AOI222_X1 port map( A1 => n3668, A2 => n8975, B1 => n6592, B2 => 
                           n8972, C1 => n3860, C2 => n8969, ZN => n1269);
   U1338 : OAI221_X1 port map( B1 => n6897, B2 => n8981, C1 => n6705, C2 => 
                           n8978, A => n2311, ZN => n2304);
   U1339 : AOI222_X1 port map( A1 => n3669, A2 => n8975, B1 => n6593, B2 => 
                           n8972, C1 => n3861, C2 => n8969, ZN => n2311);
   U1340 : OAI221_X1 port map( B1 => n6898, B2 => n8981, C1 => n6706, C2 => 
                           n8978, A => n2329, ZN => n2322);
   U1341 : AOI222_X1 port map( A1 => n3670, A2 => n8975, B1 => n6594, B2 => 
                           n8972, C1 => n3862, C2 => n8969, ZN => n2329);
   U1342 : OAI221_X1 port map( B1 => n6859, B2 => n8981, C1 => n6667, C2 => 
                           n8978, A => n2347, ZN => n2340);
   U1343 : AOI222_X1 port map( A1 => n3575, A2 => n8975, B1 => n6595, B2 => 
                           n8972, C1 => n3615, C2 => n8969, ZN => n2347);
   U1344 : OAI221_X1 port map( B1 => n6860, B2 => n8981, C1 => n6668, C2 => 
                           n8978, A => n2365, ZN => n2358);
   U1345 : AOI222_X1 port map( A1 => n3576, A2 => n8975, B1 => n6596, B2 => 
                           n8972, C1 => n3616, C2 => n8969, ZN => n2365);
   U1346 : OAI221_X1 port map( B1 => n6861, B2 => n8981, C1 => n6669, C2 => 
                           n8978, A => n2383, ZN => n2376);
   U1347 : AOI222_X1 port map( A1 => n3577, A2 => n8975, B1 => n6597, B2 => 
                           n8972, C1 => n3617, C2 => n8969, ZN => n2383);
   U1348 : OAI221_X1 port map( B1 => n6862, B2 => n8981, C1 => n6670, C2 => 
                           n8978, A => n2401, ZN => n2394);
   U1349 : AOI222_X1 port map( A1 => n3578, A2 => n8975, B1 => n6598, B2 => 
                           n8972, C1 => n3618, C2 => n8969, ZN => n2401);
   U1350 : OAI221_X1 port map( B1 => n6863, B2 => n8981, C1 => n6671, C2 => 
                           n8978, A => n2419, ZN => n2412);
   U1351 : AOI222_X1 port map( A1 => n3579, A2 => n8975, B1 => n6599, B2 => 
                           n8972, C1 => n3619, C2 => n8969, ZN => n2419);
   U1352 : OAI221_X1 port map( B1 => n6864, B2 => n8981, C1 => n6672, C2 => 
                           n8978, A => n2437, ZN => n2430);
   U1353 : AOI222_X1 port map( A1 => n3580, A2 => n8975, B1 => n6600, B2 => 
                           n8972, C1 => n3620, C2 => n8969, ZN => n2437);
   U1354 : OAI221_X1 port map( B1 => n6865, B2 => n8981, C1 => n6673, C2 => 
                           n8978, A => n2455, ZN => n2448);
   U1355 : AOI222_X1 port map( A1 => n3581, A2 => n8975, B1 => n6601, B2 => 
                           n8972, C1 => n3621, C2 => n8969, ZN => n2455);
   U1356 : OAI221_X1 port map( B1 => n6866, B2 => n8981, C1 => n6674, C2 => 
                           n8978, A => n2483, ZN => n2466);
   U1357 : AOI222_X1 port map( A1 => n3582, A2 => n8975, B1 => n6602, B2 => 
                           n8972, C1 => n3622, C2 => n8969, ZN => n2483);
   U1358 : NOR4_X1 port map( A1 => n2675, A2 => n2676, A3 => n2677, A4 => n2678
                           , ZN => n2674);
   U1359 : OAI221_X1 port map( B1 => n7798, B2 => n8883, C1 => n8037, C2 => 
                           n8880, A => n2682, ZN => n2675);
   U1360 : OAI221_X1 port map( B1 => n7797, B2 => n8895, C1 => n8005, C2 => 
                           n8892, A => n2681, ZN => n2676);
   U1361 : OAI221_X1 port map( B1 => n7981, B2 => n8919, C1 => n6755, C2 => 
                           n8916, A => n2679, ZN => n2678);
   U1362 : NOR4_X1 port map( A1 => n2693, A2 => n2694, A3 => n2695, A4 => n2696
                           , ZN => n2692);
   U1363 : OAI221_X1 port map( B1 => n7800, B2 => n8883, C1 => n8038, C2 => 
                           n8880, A => n2700, ZN => n2693);
   U1364 : OAI221_X1 port map( B1 => n7799, B2 => n8895, C1 => n8006, C2 => 
                           n8892, A => n2699, ZN => n2694);
   U1365 : OAI221_X1 port map( B1 => n7982, B2 => n8919, C1 => n6756, C2 => 
                           n8916, A => n2697, ZN => n2696);
   U1366 : NOR4_X1 port map( A1 => n2711, A2 => n2712, A3 => n2713, A4 => n2714
                           , ZN => n2710);
   U1367 : OAI221_X1 port map( B1 => n7802, B2 => n8883, C1 => n8039, C2 => 
                           n8880, A => n2718, ZN => n2711);
   U1368 : OAI221_X1 port map( B1 => n7801, B2 => n8895, C1 => n8007, C2 => 
                           n8892, A => n2717, ZN => n2712);
   U1369 : OAI221_X1 port map( B1 => n7983, B2 => n8919, C1 => n6757, C2 => 
                           n8916, A => n2715, ZN => n2714);
   U1370 : NOR4_X1 port map( A1 => n2729, A2 => n2730, A3 => n2731, A4 => n2732
                           , ZN => n2728);
   U1371 : OAI221_X1 port map( B1 => n7804, B2 => n8883, C1 => n8040, C2 => 
                           n8880, A => n2736, ZN => n2729);
   U1372 : OAI221_X1 port map( B1 => n7803, B2 => n8895, C1 => n8008, C2 => 
                           n8892, A => n2735, ZN => n2730);
   U1373 : OAI221_X1 port map( B1 => n7984, B2 => n8919, C1 => n6758, C2 => 
                           n8916, A => n2733, ZN => n2732);
   U1374 : NOR4_X1 port map( A1 => n2747, A2 => n2748, A3 => n2749, A4 => n2750
                           , ZN => n2746);
   U1375 : OAI221_X1 port map( B1 => n7658, B2 => n8883, C1 => n8041, C2 => 
                           n8880, A => n2754, ZN => n2747);
   U1376 : OAI221_X1 port map( B1 => n7657, B2 => n8895, C1 => n8009, C2 => 
                           n8892, A => n2753, ZN => n2748);
   U1377 : OAI221_X1 port map( B1 => n7985, B2 => n8919, C1 => n6759, C2 => 
                           n8916, A => n2751, ZN => n2750);
   U1378 : NOR4_X1 port map( A1 => n2765, A2 => n2766, A3 => n2767, A4 => n2768
                           , ZN => n2764);
   U1379 : OAI221_X1 port map( B1 => n7660, B2 => n8883, C1 => n8042, C2 => 
                           n8880, A => n2772, ZN => n2765);
   U1380 : OAI221_X1 port map( B1 => n7659, B2 => n8895, C1 => n8010, C2 => 
                           n8892, A => n2771, ZN => n2766);
   U1381 : OAI221_X1 port map( B1 => n7986, B2 => n8919, C1 => n6760, C2 => 
                           n8916, A => n2769, ZN => n2768);
   U1382 : NOR4_X1 port map( A1 => n2783, A2 => n2784, A3 => n2785, A4 => n2786
                           , ZN => n2782);
   U1383 : OAI221_X1 port map( B1 => n7662, B2 => n8883, C1 => n8043, C2 => 
                           n8880, A => n2790, ZN => n2783);
   U1384 : OAI221_X1 port map( B1 => n7661, B2 => n8895, C1 => n8011, C2 => 
                           n8892, A => n2789, ZN => n2784);
   U1385 : OAI221_X1 port map( B1 => n7987, B2 => n8919, C1 => n6761, C2 => 
                           n8916, A => n2787, ZN => n2786);
   U1386 : NOR4_X1 port map( A1 => n2801, A2 => n2802, A3 => n2803, A4 => n2804
                           , ZN => n2800);
   U1387 : OAI221_X1 port map( B1 => n7664, B2 => n8883, C1 => n8044, C2 => 
                           n8880, A => n2808, ZN => n2801);
   U1388 : OAI221_X1 port map( B1 => n7663, B2 => n8895, C1 => n8012, C2 => 
                           n8892, A => n2807, ZN => n2802);
   U1389 : OAI221_X1 port map( B1 => n7988, B2 => n8919, C1 => n6762, C2 => 
                           n8916, A => n2805, ZN => n2804);
   U1390 : NOR4_X1 port map( A1 => n2819, A2 => n2820, A3 => n2821, A4 => n2822
                           , ZN => n2818);
   U1391 : OAI221_X1 port map( B1 => n7666, B2 => n8883, C1 => n8045, C2 => 
                           n8880, A => n2826, ZN => n2819);
   U1392 : OAI221_X1 port map( B1 => n7665, B2 => n8895, C1 => n8013, C2 => 
                           n8892, A => n2825, ZN => n2820);
   U1393 : OAI221_X1 port map( B1 => n7989, B2 => n8919, C1 => n6763, C2 => 
                           n8916, A => n2823, ZN => n2822);
   U1394 : NOR4_X1 port map( A1 => n2837, A2 => n2838, A3 => n2839, A4 => n2840
                           , ZN => n2836);
   U1395 : OAI221_X1 port map( B1 => n7668, B2 => n8883, C1 => n8046, C2 => 
                           n8880, A => n2844, ZN => n2837);
   U1396 : OAI221_X1 port map( B1 => n7667, B2 => n8895, C1 => n8014, C2 => 
                           n8892, A => n2843, ZN => n2838);
   U1397 : OAI221_X1 port map( B1 => n7990, B2 => n8919, C1 => n6764, C2 => 
                           n8916, A => n2841, ZN => n2840);
   U1398 : NOR4_X1 port map( A1 => n2855, A2 => n2856, A3 => n2857, A4 => n2858
                           , ZN => n2854);
   U1399 : OAI221_X1 port map( B1 => n7670, B2 => n8883, C1 => n8047, C2 => 
                           n8880, A => n2862, ZN => n2855);
   U1400 : OAI221_X1 port map( B1 => n7669, B2 => n8895, C1 => n8015, C2 => 
                           n8892, A => n2861, ZN => n2856);
   U1401 : OAI221_X1 port map( B1 => n7991, B2 => n8919, C1 => n6765, C2 => 
                           n8916, A => n2859, ZN => n2858);
   U1402 : NOR4_X1 port map( A1 => n2873, A2 => n2874, A3 => n2875, A4 => n2876
                           , ZN => n2872);
   U1403 : OAI221_X1 port map( B1 => n7672, B2 => n8883, C1 => n8048, C2 => 
                           n8880, A => n2880, ZN => n2873);
   U1404 : OAI221_X1 port map( B1 => n7671, B2 => n8895, C1 => n8016, C2 => 
                           n8892, A => n2879, ZN => n2874);
   U1405 : OAI221_X1 port map( B1 => n7992, B2 => n8919, C1 => n6766, C2 => 
                           n8916, A => n2877, ZN => n2876);
   U1406 : NOR4_X1 port map( A1 => n2891, A2 => n2892, A3 => n2893, A4 => n2894
                           , ZN => n2890);
   U1407 : OAI221_X1 port map( B1 => n7674, B2 => n8882, C1 => n8049, C2 => 
                           n8879, A => n2898, ZN => n2891);
   U1408 : OAI221_X1 port map( B1 => n7673, B2 => n8894, C1 => n8017, C2 => 
                           n8891, A => n2897, ZN => n2892);
   U1409 : OAI221_X1 port map( B1 => n7993, B2 => n8918, C1 => n6767, C2 => 
                           n8915, A => n2895, ZN => n2894);
   U1410 : NOR4_X1 port map( A1 => n2909, A2 => n2910, A3 => n2911, A4 => n2912
                           , ZN => n2908);
   U1411 : OAI221_X1 port map( B1 => n7676, B2 => n8882, C1 => n8050, C2 => 
                           n8879, A => n2916, ZN => n2909);
   U1412 : OAI221_X1 port map( B1 => n7675, B2 => n8894, C1 => n8018, C2 => 
                           n8891, A => n2915, ZN => n2910);
   U1413 : OAI221_X1 port map( B1 => n7994, B2 => n8918, C1 => n6768, C2 => 
                           n8915, A => n2913, ZN => n2912);
   U1414 : NOR4_X1 port map( A1 => n2927, A2 => n2928, A3 => n2929, A4 => n2930
                           , ZN => n2926);
   U1415 : OAI221_X1 port map( B1 => n7678, B2 => n8882, C1 => n8051, C2 => 
                           n8879, A => n2934, ZN => n2927);
   U1416 : OAI221_X1 port map( B1 => n7677, B2 => n8894, C1 => n8019, C2 => 
                           n8891, A => n2933, ZN => n2928);
   U1417 : OAI221_X1 port map( B1 => n7995, B2 => n8918, C1 => n6769, C2 => 
                           n8915, A => n2931, ZN => n2930);
   U1418 : NOR4_X1 port map( A1 => n2945, A2 => n2946, A3 => n2947, A4 => n2948
                           , ZN => n2944);
   U1419 : OAI221_X1 port map( B1 => n7680, B2 => n8882, C1 => n8052, C2 => 
                           n8879, A => n2952, ZN => n2945);
   U1420 : OAI221_X1 port map( B1 => n7679, B2 => n8894, C1 => n8020, C2 => 
                           n8891, A => n2951, ZN => n2946);
   U1421 : OAI221_X1 port map( B1 => n7996, B2 => n8918, C1 => n6770, C2 => 
                           n8915, A => n2949, ZN => n2948);
   U1422 : NOR4_X1 port map( A1 => n2963, A2 => n2964, A3 => n2965, A4 => n2966
                           , ZN => n2962);
   U1423 : OAI221_X1 port map( B1 => n7681, B2 => n8882, C1 => n7821, C2 => 
                           n8879, A => n2970, ZN => n2963);
   U1424 : OAI221_X1 port map( B1 => n7806, B2 => n8894, C1 => n8021, C2 => 
                           n8891, A => n2969, ZN => n2964);
   U1425 : OAI221_X1 port map( B1 => n7805, B2 => n8918, C1 => n6731, C2 => 
                           n8915, A => n2967, ZN => n2966);
   U1426 : NOR4_X1 port map( A1 => n2981, A2 => n2982, A3 => n2983, A4 => n2984
                           , ZN => n2980);
   U1427 : OAI221_X1 port map( B1 => n7682, B2 => n8882, C1 => n7822, C2 => 
                           n8879, A => n2988, ZN => n2981);
   U1428 : OAI221_X1 port map( B1 => n7808, B2 => n8894, C1 => n8022, C2 => 
                           n8891, A => n2987, ZN => n2982);
   U1429 : OAI221_X1 port map( B1 => n7807, B2 => n8918, C1 => n6732, C2 => 
                           n8915, A => n2985, ZN => n2984);
   U1430 : NOR4_X1 port map( A1 => n2999, A2 => n3000, A3 => n3001, A4 => n3002
                           , ZN => n2998);
   U1431 : OAI221_X1 port map( B1 => n7683, B2 => n8882, C1 => n7823, C2 => 
                           n8879, A => n3006, ZN => n2999);
   U1432 : OAI221_X1 port map( B1 => n7810, B2 => n8894, C1 => n8023, C2 => 
                           n8891, A => n3005, ZN => n3000);
   U1433 : OAI221_X1 port map( B1 => n7809, B2 => n8918, C1 => n6733, C2 => 
                           n8915, A => n3003, ZN => n3002);
   U1434 : NOR4_X1 port map( A1 => n3017, A2 => n3018, A3 => n3019, A4 => n3020
                           , ZN => n3016);
   U1435 : OAI221_X1 port map( B1 => n7684, B2 => n8882, C1 => n7824, C2 => 
                           n8879, A => n3024, ZN => n3017);
   U1436 : OAI221_X1 port map( B1 => n7812, B2 => n8894, C1 => n8024, C2 => 
                           n8891, A => n3023, ZN => n3018);
   U1437 : OAI221_X1 port map( B1 => n7811, B2 => n8918, C1 => n6734, C2 => 
                           n8915, A => n3021, ZN => n3020);
   U1438 : NOR4_X1 port map( A1 => n3035, A2 => n3036, A3 => n3037, A4 => n3038
                           , ZN => n3034);
   U1439 : OAI221_X1 port map( B1 => n7685, B2 => n8882, C1 => n7825, C2 => 
                           n8879, A => n3042, ZN => n3035);
   U1440 : OAI221_X1 port map( B1 => n7814, B2 => n8894, C1 => n8025, C2 => 
                           n8891, A => n3041, ZN => n3036);
   U1441 : OAI221_X1 port map( B1 => n7813, B2 => n8918, C1 => n6735, C2 => 
                           n8915, A => n3039, ZN => n3038);
   U1442 : NOR4_X1 port map( A1 => n3053, A2 => n3054, A3 => n3055, A4 => n3056
                           , ZN => n3052);
   U1443 : OAI221_X1 port map( B1 => n7686, B2 => n8882, C1 => n7826, C2 => 
                           n8879, A => n3060, ZN => n3053);
   U1444 : OAI221_X1 port map( B1 => n7816, B2 => n8894, C1 => n8026, C2 => 
                           n8891, A => n3059, ZN => n3054);
   U1445 : OAI221_X1 port map( B1 => n7815, B2 => n8918, C1 => n6736, C2 => 
                           n8915, A => n3057, ZN => n3056);
   U1446 : NOR4_X1 port map( A1 => n3071, A2 => n3072, A3 => n3073, A4 => n3074
                           , ZN => n3070);
   U1447 : OAI221_X1 port map( B1 => n7687, B2 => n8882, C1 => n7827, C2 => 
                           n8879, A => n3078, ZN => n3071);
   U1448 : OAI221_X1 port map( B1 => n7818, B2 => n8894, C1 => n8027, C2 => 
                           n8891, A => n3077, ZN => n3072);
   U1449 : OAI221_X1 port map( B1 => n7817, B2 => n8918, C1 => n6737, C2 => 
                           n8915, A => n3075, ZN => n3074);
   U1450 : NOR4_X1 port map( A1 => n3089, A2 => n3090, A3 => n3091, A4 => n3092
                           , ZN => n3088);
   U1451 : OAI221_X1 port map( B1 => n7688, B2 => n8882, C1 => n7828, C2 => 
                           n8879, A => n3104, ZN => n3089);
   U1452 : OAI221_X1 port map( B1 => n7820, B2 => n8894, C1 => n8028, C2 => 
                           n8891, A => n3101, ZN => n3090);
   U1453 : OAI221_X1 port map( B1 => n7819, B2 => n8918, C1 => n6738, C2 => 
                           n8915, A => n3093, ZN => n3092);
   U1454 : NOR4_X1 port map( A1 => n2498, A2 => n2499, A3 => n2500, A4 => n2501
                           , ZN => n2497);
   U1455 : OAI221_X1 port map( B1 => n7781, B2 => n8884, C1 => n8029, C2 => 
                           n8881, A => n2519, ZN => n2498);
   U1456 : OAI221_X1 port map( B1 => n7789, B2 => n8896, C1 => n7997, C2 => 
                           n8893, A => n2514, ZN => n2499);
   U1457 : OAI221_X1 port map( B1 => n7973, B2 => n8920, C1 => n6747, C2 => 
                           n8917, A => n2504, ZN => n2501);
   U1458 : NOR4_X1 port map( A1 => n2549, A2 => n2550, A3 => n2551, A4 => n2552
                           , ZN => n2548);
   U1459 : OAI221_X1 port map( B1 => n7782, B2 => n8884, C1 => n8030, C2 => 
                           n8881, A => n2556, ZN => n2549);
   U1460 : OAI221_X1 port map( B1 => n7790, B2 => n8896, C1 => n7998, C2 => 
                           n8893, A => n2555, ZN => n2550);
   U1461 : OAI221_X1 port map( B1 => n7974, B2 => n8920, C1 => n6748, C2 => 
                           n8917, A => n2553, ZN => n2552);
   U1462 : NOR4_X1 port map( A1 => n2567, A2 => n2568, A3 => n2569, A4 => n2570
                           , ZN => n2566);
   U1463 : OAI221_X1 port map( B1 => n7783, B2 => n8884, C1 => n8031, C2 => 
                           n8881, A => n2574, ZN => n2567);
   U1464 : OAI221_X1 port map( B1 => n7791, B2 => n8896, C1 => n7999, C2 => 
                           n8893, A => n2573, ZN => n2568);
   U1465 : OAI221_X1 port map( B1 => n7975, B2 => n8920, C1 => n6749, C2 => 
                           n8917, A => n2571, ZN => n2570);
   U1466 : NOR4_X1 port map( A1 => n2585, A2 => n2586, A3 => n2587, A4 => n2588
                           , ZN => n2584);
   U1467 : OAI221_X1 port map( B1 => n7784, B2 => n8884, C1 => n8032, C2 => 
                           n8881, A => n2592, ZN => n2585);
   U1468 : OAI221_X1 port map( B1 => n7792, B2 => n8896, C1 => n8000, C2 => 
                           n8893, A => n2591, ZN => n2586);
   U1469 : OAI221_X1 port map( B1 => n7976, B2 => n8920, C1 => n6750, C2 => 
                           n8917, A => n2589, ZN => n2588);
   U1470 : NOR4_X1 port map( A1 => n2603, A2 => n2604, A3 => n2605, A4 => n2606
                           , ZN => n2602);
   U1471 : OAI221_X1 port map( B1 => n7785, B2 => n8884, C1 => n8033, C2 => 
                           n8881, A => n2610, ZN => n2603);
   U1472 : OAI221_X1 port map( B1 => n7793, B2 => n8896, C1 => n8001, C2 => 
                           n8893, A => n2609, ZN => n2604);
   U1473 : OAI221_X1 port map( B1 => n7977, B2 => n8920, C1 => n6751, C2 => 
                           n8917, A => n2607, ZN => n2606);
   U1474 : NOR4_X1 port map( A1 => n2621, A2 => n2622, A3 => n2623, A4 => n2624
                           , ZN => n2620);
   U1475 : OAI221_X1 port map( B1 => n7786, B2 => n8884, C1 => n8034, C2 => 
                           n8881, A => n2628, ZN => n2621);
   U1476 : OAI221_X1 port map( B1 => n7794, B2 => n8896, C1 => n8002, C2 => 
                           n8893, A => n2627, ZN => n2622);
   U1477 : OAI221_X1 port map( B1 => n7978, B2 => n8920, C1 => n6752, C2 => 
                           n8917, A => n2625, ZN => n2624);
   U1478 : NOR4_X1 port map( A1 => n2639, A2 => n2640, A3 => n2641, A4 => n2642
                           , ZN => n2638);
   U1479 : OAI221_X1 port map( B1 => n7787, B2 => n8884, C1 => n8035, C2 => 
                           n8881, A => n2646, ZN => n2639);
   U1480 : OAI221_X1 port map( B1 => n7795, B2 => n8896, C1 => n8003, C2 => 
                           n8893, A => n2645, ZN => n2640);
   U1481 : OAI221_X1 port map( B1 => n7979, B2 => n8920, C1 => n6753, C2 => 
                           n8917, A => n2643, ZN => n2642);
   U1482 : NOR4_X1 port map( A1 => n2657, A2 => n2658, A3 => n2659, A4 => n2660
                           , ZN => n2656);
   U1483 : OAI221_X1 port map( B1 => n7788, B2 => n8884, C1 => n8036, C2 => 
                           n8881, A => n2664, ZN => n2657);
   U1484 : OAI221_X1 port map( B1 => n7796, B2 => n8896, C1 => n8004, C2 => 
                           n8893, A => n2663, ZN => n2658);
   U1485 : OAI221_X1 port map( B1 => n7980, B2 => n8920, C1 => n6754, C2 => 
                           n8917, A => n2661, ZN => n2660);
   U1486 : OAI221_X1 port map( B1 => n8956, B2 => n8133, C1 => n6771, C2 => 
                           n8953, A => n887, ZN => n878);
   U1487 : AOI22_X1 port map( A1 => n8950, A2 => n8229, B1 => n3311, B2 => 
                           n8947, ZN => n887);
   U1488 : OAI221_X1 port map( B1 => n8956, B2 => n8134, C1 => n6772, C2 => 
                           n8953, A => n915, ZN => n912);
   U1489 : AOI22_X1 port map( A1 => n8950, A2 => n8230, B1 => n3312, B2 => 
                           n8947, ZN => n915);
   U1490 : OAI221_X1 port map( B1 => n8956, B2 => n8135, C1 => n6773, C2 => 
                           n8953, A => n933, ZN => n930);
   U1491 : AOI22_X1 port map( A1 => n8950, A2 => n8231, B1 => n3313, B2 => 
                           n8947, ZN => n933);
   U1492 : OAI221_X1 port map( B1 => n8956, B2 => n8136, C1 => n6774, C2 => 
                           n8953, A => n951, ZN => n948);
   U1493 : AOI22_X1 port map( A1 => n8950, A2 => n8232, B1 => n3314, B2 => 
                           n8947, ZN => n951);
   U1494 : OAI221_X1 port map( B1 => n8956, B2 => n8137, C1 => n6775, C2 => 
                           n8953, A => n969, ZN => n966);
   U1495 : AOI22_X1 port map( A1 => n8950, A2 => n8233, B1 => n3315, B2 => 
                           n8947, ZN => n969);
   U1496 : OAI221_X1 port map( B1 => n8956, B2 => n8138, C1 => n6776, C2 => 
                           n8953, A => n987, ZN => n984);
   U1497 : AOI22_X1 port map( A1 => n8950, A2 => n8234, B1 => n3316, B2 => 
                           n8947, ZN => n987);
   U1498 : OAI221_X1 port map( B1 => n8956, B2 => n8139, C1 => n6777, C2 => 
                           n8953, A => n1005, ZN => n1002);
   U1499 : AOI22_X1 port map( A1 => n8950, A2 => n8235, B1 => n3317, B2 => 
                           n8947, ZN => n1005);
   U1500 : OAI221_X1 port map( B1 => n8956, B2 => n8140, C1 => n6778, C2 => 
                           n8953, A => n1023, ZN => n1020);
   U1501 : AOI22_X1 port map( A1 => n8950, A2 => n8236, B1 => n3318, B2 => 
                           n8947, ZN => n1023);
   U1502 : OAI221_X1 port map( B1 => n6627, B2 => n9007, C1 => n6339, C2 => 
                           n9004, A => n862, ZN => n853);
   U1503 : AOI22_X1 port map( A1 => n3719, A2 => n9001, B1 => n3623, B2 => 
                           n8998, ZN => n862);
   U1504 : OAI221_X1 port map( B1 => n6628, B2 => n9007, C1 => n6340, C2 => 
                           n9004, A => n907, ZN => n904);
   U1505 : AOI22_X1 port map( A1 => n3720, A2 => n9001, B1 => n3624, B2 => 
                           n8998, ZN => n907);
   U1506 : OAI221_X1 port map( B1 => n6629, B2 => n9007, C1 => n6341, C2 => 
                           n9004, A => n925, ZN => n922);
   U1507 : AOI22_X1 port map( A1 => n3721, A2 => n9001, B1 => n3625, B2 => 
                           n8998, ZN => n925);
   U1508 : OAI221_X1 port map( B1 => n6630, B2 => n9007, C1 => n6342, C2 => 
                           n9004, A => n943, ZN => n940);
   U1509 : AOI22_X1 port map( A1 => n3722, A2 => n9001, B1 => n3626, B2 => 
                           n8998, ZN => n943);
   U1510 : OAI221_X1 port map( B1 => n6631, B2 => n9007, C1 => n6343, C2 => 
                           n9004, A => n961, ZN => n958);
   U1511 : AOI22_X1 port map( A1 => n3723, A2 => n9001, B1 => n3627, B2 => 
                           n8998, ZN => n961);
   U1512 : OAI221_X1 port map( B1 => n6632, B2 => n9007, C1 => n6344, C2 => 
                           n9004, A => n979, ZN => n976);
   U1513 : AOI22_X1 port map( A1 => n3724, A2 => n9001, B1 => n3628, B2 => 
                           n8998, ZN => n979);
   U1514 : OAI221_X1 port map( B1 => n6633, B2 => n9007, C1 => n6345, C2 => 
                           n9004, A => n997, ZN => n994);
   U1515 : AOI22_X1 port map( A1 => n3725, A2 => n9001, B1 => n3629, B2 => 
                           n8998, ZN => n997);
   U1516 : OAI221_X1 port map( B1 => n6634, B2 => n9007, C1 => n6346, C2 => 
                           n9004, A => n1015, ZN => n1012);
   U1517 : AOI22_X1 port map( A1 => n3726, A2 => n9001, B1 => n3630, B2 => 
                           n8998, ZN => n1015);
   U1518 : OAI221_X1 port map( B1 => n6603, B2 => n9006, C1 => n6315, C2 => 
                           n9003, A => n1033, ZN => n1030);
   U1519 : AOI22_X1 port map( A1 => n3727, A2 => n9000, B1 => n3631, B2 => 
                           n8997, ZN => n1033);
   U1520 : OAI221_X1 port map( B1 => n6604, B2 => n9006, C1 => n6316, C2 => 
                           n9003, A => n1051, ZN => n1048);
   U1521 : AOI22_X1 port map( A1 => n3728, A2 => n9000, B1 => n3632, B2 => 
                           n8997, ZN => n1051);
   U1522 : OAI221_X1 port map( B1 => n6605, B2 => n9006, C1 => n6317, C2 => 
                           n9003, A => n1069, ZN => n1066);
   U1523 : AOI22_X1 port map( A1 => n3729, A2 => n9000, B1 => n3633, B2 => 
                           n8997, ZN => n1069);
   U1524 : OAI221_X1 port map( B1 => n6606, B2 => n9006, C1 => n6318, C2 => 
                           n9003, A => n1087, ZN => n1084);
   U1525 : AOI22_X1 port map( A1 => n3730, A2 => n9000, B1 => n3634, B2 => 
                           n8997, ZN => n1087);
   U1526 : OAI221_X1 port map( B1 => n6607, B2 => n9006, C1 => n6319, C2 => 
                           n9003, A => n1105, ZN => n1102);
   U1527 : AOI22_X1 port map( A1 => n3731, A2 => n9000, B1 => n3635, B2 => 
                           n8997, ZN => n1105);
   U1528 : OAI221_X1 port map( B1 => n6608, B2 => n9006, C1 => n6320, C2 => 
                           n9003, A => n1123, ZN => n1120);
   U1529 : AOI22_X1 port map( A1 => n3732, A2 => n9000, B1 => n3636, B2 => 
                           n8997, ZN => n1123);
   U1530 : OAI221_X1 port map( B1 => n6609, B2 => n9006, C1 => n6321, C2 => 
                           n9003, A => n1141, ZN => n1138);
   U1531 : AOI22_X1 port map( A1 => n3733, A2 => n9000, B1 => n3637, B2 => 
                           n8997, ZN => n1141);
   U1532 : OAI221_X1 port map( B1 => n6610, B2 => n9006, C1 => n6322, C2 => 
                           n9003, A => n1159, ZN => n1156);
   U1533 : AOI22_X1 port map( A1 => n3734, A2 => n9000, B1 => n3638, B2 => 
                           n8997, ZN => n1159);
   U1534 : OAI221_X1 port map( B1 => n6611, B2 => n9006, C1 => n6323, C2 => 
                           n9003, A => n1177, ZN => n1174);
   U1535 : AOI22_X1 port map( A1 => n3735, A2 => n9000, B1 => n3639, B2 => 
                           n8997, ZN => n1177);
   U1536 : OAI221_X1 port map( B1 => n6612, B2 => n9006, C1 => n6324, C2 => 
                           n9003, A => n1195, ZN => n1192);
   U1537 : AOI22_X1 port map( A1 => n3736, A2 => n9000, B1 => n3640, B2 => 
                           n8997, ZN => n1195);
   U1538 : OAI221_X1 port map( B1 => n6613, B2 => n9006, C1 => n6325, C2 => 
                           n9003, A => n1213, ZN => n1210);
   U1539 : AOI22_X1 port map( A1 => n3737, A2 => n9000, B1 => n3641, B2 => 
                           n8997, ZN => n1213);
   U1540 : OAI221_X1 port map( B1 => n6614, B2 => n9006, C1 => n6326, C2 => 
                           n9003, A => n1231, ZN => n1228);
   U1541 : AOI22_X1 port map( A1 => n3738, A2 => n9000, B1 => n3642, B2 => 
                           n8997, ZN => n1231);
   U1542 : OAI221_X1 port map( B1 => n6615, B2 => n9005, C1 => n6327, C2 => 
                           n9002, A => n1249, ZN => n1246);
   U1543 : AOI22_X1 port map( A1 => n3739, A2 => n8999, B1 => n3643, B2 => 
                           n8996, ZN => n1249);
   U1544 : OAI221_X1 port map( B1 => n6616, B2 => n9005, C1 => n6328, C2 => 
                           n9002, A => n1267, ZN => n1264);
   U1545 : AOI22_X1 port map( A1 => n3740, A2 => n8999, B1 => n3644, B2 => 
                           n8996, ZN => n1267);
   U1546 : OAI221_X1 port map( B1 => n6617, B2 => n9005, C1 => n6329, C2 => 
                           n9002, A => n2309, ZN => n2306);
   U1547 : AOI22_X1 port map( A1 => n3741, A2 => n8999, B1 => n3645, B2 => 
                           n8996, ZN => n2309);
   U1548 : OAI221_X1 port map( B1 => n6618, B2 => n9005, C1 => n6330, C2 => 
                           n9002, A => n2327, ZN => n2324);
   U1549 : AOI22_X1 port map( A1 => n3742, A2 => n8999, B1 => n3646, B2 => 
                           n8996, ZN => n2327);
   U1550 : OAI221_X1 port map( B1 => n6619, B2 => n9005, C1 => n6331, C2 => 
                           n9002, A => n2345, ZN => n2342);
   U1551 : AOI22_X1 port map( A1 => n3543, A2 => n8999, B1 => n3551, B2 => 
                           n8996, ZN => n2345);
   U1552 : OAI221_X1 port map( B1 => n6620, B2 => n9005, C1 => n6332, C2 => 
                           n9002, A => n2363, ZN => n2360);
   U1553 : AOI22_X1 port map( A1 => n3544, A2 => n8999, B1 => n3552, B2 => 
                           n8996, ZN => n2363);
   U1554 : OAI221_X1 port map( B1 => n6621, B2 => n9005, C1 => n6333, C2 => 
                           n9002, A => n2381, ZN => n2378);
   U1555 : AOI22_X1 port map( A1 => n3545, A2 => n8999, B1 => n3553, B2 => 
                           n8996, ZN => n2381);
   U1556 : OAI221_X1 port map( B1 => n6622, B2 => n9005, C1 => n6334, C2 => 
                           n9002, A => n2399, ZN => n2396);
   U1557 : AOI22_X1 port map( A1 => n3546, A2 => n8999, B1 => n3554, B2 => 
                           n8996, ZN => n2399);
   U1558 : OAI221_X1 port map( B1 => n6623, B2 => n9005, C1 => n6335, C2 => 
                           n9002, A => n2417, ZN => n2414);
   U1559 : AOI22_X1 port map( A1 => n3547, A2 => n8999, B1 => n3555, B2 => 
                           n8996, ZN => n2417);
   U1560 : OAI221_X1 port map( B1 => n6624, B2 => n9005, C1 => n6336, C2 => 
                           n9002, A => n2435, ZN => n2432);
   U1561 : AOI22_X1 port map( A1 => n3548, A2 => n8999, B1 => n3556, B2 => 
                           n8996, ZN => n2435);
   U1562 : OAI221_X1 port map( B1 => n6625, B2 => n9005, C1 => n6337, C2 => 
                           n9002, A => n2453, ZN => n2450);
   U1563 : AOI22_X1 port map( A1 => n3549, A2 => n8999, B1 => n3557, B2 => 
                           n8996, ZN => n2453);
   U1564 : OAI221_X1 port map( B1 => n6626, B2 => n9005, C1 => n6338, C2 => 
                           n9002, A => n2477, ZN => n2468);
   U1565 : AOI22_X1 port map( A1 => n3550, A2 => n8999, B1 => n3558, B2 => 
                           n8996, ZN => n2477);
   U1566 : OAI221_X1 port map( B1 => n8932, B2 => n7781, C1 => n8929, C2 => 
                           n8029, A => n897, ZN => n876);
   U1567 : AOI22_X1 port map( A1 => n3479, A2 => n8926, B1 => n3767, B2 => 
                           n8923, ZN => n897);
   U1568 : OAI221_X1 port map( B1 => n8932, B2 => n7782, C1 => n8929, C2 => 
                           n8030, A => n917, ZN => n910);
   U1569 : AOI22_X1 port map( A1 => n3480, A2 => n8926, B1 => n3768, B2 => 
                           n8923, ZN => n917);
   U1570 : OAI221_X1 port map( B1 => n8932, B2 => n7783, C1 => n8929, C2 => 
                           n8031, A => n935, ZN => n928);
   U1571 : AOI22_X1 port map( A1 => n3481, A2 => n8926, B1 => n3769, B2 => 
                           n8923, ZN => n935);
   U1572 : OAI221_X1 port map( B1 => n8932, B2 => n7784, C1 => n8929, C2 => 
                           n8032, A => n953, ZN => n946);
   U1573 : AOI22_X1 port map( A1 => n3482, A2 => n8926, B1 => n3770, B2 => 
                           n8923, ZN => n953);
   U1574 : OAI221_X1 port map( B1 => n8932, B2 => n7785, C1 => n8929, C2 => 
                           n8033, A => n971, ZN => n964);
   U1575 : AOI22_X1 port map( A1 => n3483, A2 => n8926, B1 => n3771, B2 => 
                           n8923, ZN => n971);
   U1576 : OAI221_X1 port map( B1 => n8932, B2 => n7786, C1 => n8929, C2 => 
                           n8034, A => n989, ZN => n982);
   U1577 : AOI22_X1 port map( A1 => n3484, A2 => n8926, B1 => n3772, B2 => 
                           n8923, ZN => n989);
   U1578 : OAI221_X1 port map( B1 => n8932, B2 => n7787, C1 => n8929, C2 => 
                           n8035, A => n1007, ZN => n1000);
   U1579 : AOI22_X1 port map( A1 => n3485, A2 => n8926, B1 => n3773, B2 => 
                           n8923, ZN => n1007);
   U1580 : OAI221_X1 port map( B1 => n8932, B2 => n7788, C1 => n8929, C2 => 
                           n8036, A => n1025, ZN => n1018);
   U1581 : AOI22_X1 port map( A1 => n3486, A2 => n8926, B1 => n3774, B2 => 
                           n8923, ZN => n1025);
   U1582 : OAI221_X1 port map( B1 => n6875, B2 => n8983, C1 => n6683, C2 => 
                           n8980, A => n872, ZN => n851);
   U1583 : AOI222_X1 port map( A1 => n3647, A2 => n8977, B1 => n6571, B2 => 
                           n8974, C1 => n3839, C2 => n8971, ZN => n872);
   U1584 : OAI221_X1 port map( B1 => n6876, B2 => n8983, C1 => n6684, C2 => 
                           n8980, A => n909, ZN => n902);
   U1585 : AOI222_X1 port map( A1 => n3648, A2 => n8977, B1 => n6572, B2 => 
                           n8974, C1 => n3840, C2 => n8971, ZN => n909);
   U1586 : OAI221_X1 port map( B1 => n6877, B2 => n8983, C1 => n6685, C2 => 
                           n8980, A => n927, ZN => n920);
   U1587 : AOI222_X1 port map( A1 => n3649, A2 => n8977, B1 => n6573, B2 => 
                           n8974, C1 => n3841, C2 => n8971, ZN => n927);
   U1588 : OAI221_X1 port map( B1 => n6878, B2 => n8983, C1 => n6686, C2 => 
                           n8980, A => n945, ZN => n938);
   U1589 : AOI222_X1 port map( A1 => n3650, A2 => n8977, B1 => n6574, B2 => 
                           n8974, C1 => n3842, C2 => n8971, ZN => n945);
   U1590 : OAI221_X1 port map( B1 => n6879, B2 => n8983, C1 => n6687, C2 => 
                           n8980, A => n963, ZN => n956);
   U1591 : AOI222_X1 port map( A1 => n3651, A2 => n8977, B1 => n6575, B2 => 
                           n8974, C1 => n3843, C2 => n8971, ZN => n963);
   U1592 : OAI221_X1 port map( B1 => n6880, B2 => n8983, C1 => n6688, C2 => 
                           n8980, A => n981, ZN => n974);
   U1593 : AOI222_X1 port map( A1 => n3652, A2 => n8977, B1 => n6576, B2 => 
                           n8974, C1 => n3844, C2 => n8971, ZN => n981);
   U1594 : OAI221_X1 port map( B1 => n6881, B2 => n8983, C1 => n6689, C2 => 
                           n8980, A => n999, ZN => n992);
   U1595 : AOI222_X1 port map( A1 => n3653, A2 => n8977, B1 => n6577, B2 => 
                           n8974, C1 => n3845, C2 => n8971, ZN => n999);
   U1596 : OAI221_X1 port map( B1 => n6882, B2 => n8983, C1 => n6690, C2 => 
                           n8980, A => n1017, ZN => n1010);
   U1597 : AOI222_X1 port map( A1 => n3654, A2 => n8977, B1 => n6578, B2 => 
                           n8974, C1 => n3846, C2 => n8971, ZN => n1017);
   U1598 : OAI22_X1 port map( A1 => n6707, A2 => n8872, B1 => n6899, B2 => 
                           n8869, ZN => n2525);
   U1599 : OAI22_X1 port map( A1 => n6708, A2 => n8872, B1 => n6900, B2 => 
                           n8869, ZN => n2560);
   U1600 : OAI22_X1 port map( A1 => n6709, A2 => n8872, B1 => n6901, B2 => 
                           n8869, ZN => n2578);
   U1601 : OAI22_X1 port map( A1 => n6710, A2 => n8872, B1 => n6902, B2 => 
                           n8869, ZN => n2596);
   U1602 : OAI22_X1 port map( A1 => n6711, A2 => n8872, B1 => n6903, B2 => 
                           n8869, ZN => n2614);
   U1603 : OAI22_X1 port map( A1 => n6712, A2 => n8872, B1 => n6904, B2 => 
                           n8869, ZN => n2632);
   U1604 : OAI22_X1 port map( A1 => n6713, A2 => n8872, B1 => n6905, B2 => 
                           n8869, ZN => n2650);
   U1605 : OAI22_X1 port map( A1 => n6714, A2 => n8872, B1 => n6906, B2 => 
                           n8869, ZN => n2668);
   U1606 : OAI22_X1 port map( A1 => n6715, A2 => n8871, B1 => n6907, B2 => 
                           n8868, ZN => n2686);
   U1607 : OAI22_X1 port map( A1 => n6716, A2 => n8871, B1 => n6908, B2 => 
                           n8868, ZN => n2704);
   U1608 : OAI22_X1 port map( A1 => n6717, A2 => n8871, B1 => n6909, B2 => 
                           n8868, ZN => n2722);
   U1609 : OAI22_X1 port map( A1 => n6718, A2 => n8871, B1 => n6910, B2 => 
                           n8868, ZN => n2740);
   U1610 : OAI22_X1 port map( A1 => n6719, A2 => n8871, B1 => n6911, B2 => 
                           n8868, ZN => n2758);
   U1611 : OAI22_X1 port map( A1 => n6720, A2 => n8871, B1 => n6912, B2 => 
                           n8868, ZN => n2776);
   U1612 : OAI22_X1 port map( A1 => n6721, A2 => n8871, B1 => n6913, B2 => 
                           n8868, ZN => n2794);
   U1613 : OAI22_X1 port map( A1 => n6722, A2 => n8871, B1 => n6914, B2 => 
                           n8868, ZN => n2812);
   U1614 : OAI22_X1 port map( A1 => n6723, A2 => n8871, B1 => n6915, B2 => 
                           n8868, ZN => n2830);
   U1615 : OAI22_X1 port map( A1 => n6724, A2 => n8871, B1 => n6916, B2 => 
                           n8868, ZN => n2848);
   U1616 : OAI22_X1 port map( A1 => n6725, A2 => n8871, B1 => n6917, B2 => 
                           n8868, ZN => n2866);
   U1617 : OAI22_X1 port map( A1 => n6726, A2 => n8871, B1 => n6918, B2 => 
                           n8868, ZN => n2884);
   U1618 : OAI22_X1 port map( A1 => n6727, A2 => n8870, B1 => n6919, B2 => 
                           n8867, ZN => n2902);
   U1619 : OAI22_X1 port map( A1 => n6728, A2 => n8870, B1 => n6920, B2 => 
                           n8867, ZN => n2920);
   U1620 : OAI22_X1 port map( A1 => n6729, A2 => n8870, B1 => n6921, B2 => 
                           n8867, ZN => n2938);
   U1621 : OAI22_X1 port map( A1 => n6730, A2 => n8870, B1 => n6922, B2 => 
                           n8867, ZN => n2956);
   U1622 : OAI22_X1 port map( A1 => n6675, A2 => n8870, B1 => n6867, B2 => 
                           n8867, ZN => n2974);
   U1623 : OAI22_X1 port map( A1 => n6676, A2 => n8870, B1 => n6868, B2 => 
                           n8867, ZN => n2992);
   U1624 : OAI22_X1 port map( A1 => n6677, A2 => n8870, B1 => n6869, B2 => 
                           n8867, ZN => n3010);
   U1625 : OAI22_X1 port map( A1 => n6678, A2 => n8870, B1 => n6870, B2 => 
                           n8867, ZN => n3028);
   U1626 : OAI22_X1 port map( A1 => n6679, A2 => n8870, B1 => n6871, B2 => 
                           n8867, ZN => n3046);
   U1627 : OAI22_X1 port map( A1 => n6680, A2 => n8870, B1 => n6872, B2 => 
                           n8867, ZN => n3064);
   U1628 : OAI22_X1 port map( A1 => n6681, A2 => n8870, B1 => n6873, B2 => 
                           n8867, ZN => n3082);
   U1629 : OAI22_X1 port map( A1 => n6682, A2 => n8870, B1 => n6874, B2 => 
                           n8867, ZN => n3111);
   U1630 : OAI22_X1 port map( A1 => n6339, A2 => n8827, B1 => n6627, B2 => 
                           n8824, ZN => n2542);
   U1631 : OAI22_X1 port map( A1 => n6340, A2 => n8827, B1 => n6628, B2 => 
                           n8824, ZN => n2562);
   U1632 : OAI22_X1 port map( A1 => n6341, A2 => n8827, B1 => n6629, B2 => 
                           n8824, ZN => n2580);
   U1633 : OAI22_X1 port map( A1 => n6342, A2 => n8827, B1 => n6630, B2 => 
                           n8824, ZN => n2598);
   U1634 : OAI22_X1 port map( A1 => n6343, A2 => n8827, B1 => n6631, B2 => 
                           n8824, ZN => n2616);
   U1635 : OAI22_X1 port map( A1 => n6344, A2 => n8827, B1 => n6632, B2 => 
                           n8824, ZN => n2634);
   U1636 : OAI22_X1 port map( A1 => n6345, A2 => n8827, B1 => n6633, B2 => 
                           n8824, ZN => n2652);
   U1637 : OAI22_X1 port map( A1 => n6346, A2 => n8827, B1 => n6634, B2 => 
                           n8824, ZN => n2670);
   U1638 : OAI22_X1 port map( A1 => n6315, A2 => n8826, B1 => n6603, B2 => 
                           n8823, ZN => n2688);
   U1639 : OAI22_X1 port map( A1 => n6316, A2 => n8826, B1 => n6604, B2 => 
                           n8823, ZN => n2706);
   U1640 : OAI22_X1 port map( A1 => n6317, A2 => n8826, B1 => n6605, B2 => 
                           n8823, ZN => n2724);
   U1641 : OAI22_X1 port map( A1 => n6318, A2 => n8826, B1 => n6606, B2 => 
                           n8823, ZN => n2742);
   U1642 : OAI22_X1 port map( A1 => n6319, A2 => n8826, B1 => n6607, B2 => 
                           n8823, ZN => n2760);
   U1643 : OAI22_X1 port map( A1 => n6320, A2 => n8826, B1 => n6608, B2 => 
                           n8823, ZN => n2778);
   U1644 : OAI22_X1 port map( A1 => n6321, A2 => n8826, B1 => n6609, B2 => 
                           n8823, ZN => n2796);
   U1645 : OAI22_X1 port map( A1 => n6322, A2 => n8826, B1 => n6610, B2 => 
                           n8823, ZN => n2814);
   U1646 : OAI22_X1 port map( A1 => n6323, A2 => n8826, B1 => n6611, B2 => 
                           n8823, ZN => n2832);
   U1647 : OAI22_X1 port map( A1 => n6324, A2 => n8826, B1 => n6612, B2 => 
                           n8823, ZN => n2850);
   U1648 : OAI22_X1 port map( A1 => n6325, A2 => n8826, B1 => n6613, B2 => 
                           n8823, ZN => n2868);
   U1649 : OAI22_X1 port map( A1 => n6326, A2 => n8826, B1 => n6614, B2 => 
                           n8823, ZN => n2886);
   U1650 : OAI22_X1 port map( A1 => n6327, A2 => n8825, B1 => n6615, B2 => 
                           n8822, ZN => n2904);
   U1651 : OAI22_X1 port map( A1 => n6328, A2 => n8825, B1 => n6616, B2 => 
                           n8822, ZN => n2922);
   U1652 : OAI22_X1 port map( A1 => n6329, A2 => n8825, B1 => n6617, B2 => 
                           n8822, ZN => n2940);
   U1653 : OAI22_X1 port map( A1 => n6330, A2 => n8825, B1 => n6618, B2 => 
                           n8822, ZN => n2958);
   U1654 : OAI22_X1 port map( A1 => n6331, A2 => n8825, B1 => n6619, B2 => 
                           n8822, ZN => n2976);
   U1655 : OAI22_X1 port map( A1 => n6332, A2 => n8825, B1 => n6620, B2 => 
                           n8822, ZN => n2994);
   U1656 : OAI22_X1 port map( A1 => n6333, A2 => n8825, B1 => n6621, B2 => 
                           n8822, ZN => n3012);
   U1657 : OAI22_X1 port map( A1 => n6334, A2 => n8825, B1 => n6622, B2 => 
                           n8822, ZN => n3030);
   U1658 : OAI22_X1 port map( A1 => n6335, A2 => n8825, B1 => n6623, B2 => 
                           n8822, ZN => n3048);
   U1659 : OAI22_X1 port map( A1 => n6336, A2 => n8825, B1 => n6624, B2 => 
                           n8822, ZN => n3066);
   U1660 : OAI22_X1 port map( A1 => n6337, A2 => n8825, B1 => n6625, B2 => 
                           n8822, ZN => n3084);
   U1661 : OAI22_X1 port map( A1 => n6338, A2 => n8825, B1 => n6626, B2 => 
                           n8822, ZN => n3114);
   U1662 : OAI22_X1 port map( A1 => n6683, A2 => n8860, B1 => n6875, B2 => 
                           n8857, ZN => n2523);
   U1663 : OAI22_X1 port map( A1 => n6684, A2 => n8860, B1 => n6876, B2 => 
                           n8857, ZN => n2558);
   U1664 : OAI22_X1 port map( A1 => n6685, A2 => n8860, B1 => n6877, B2 => 
                           n8857, ZN => n2576);
   U1665 : OAI22_X1 port map( A1 => n6686, A2 => n8860, B1 => n6878, B2 => 
                           n8857, ZN => n2594);
   U1666 : OAI22_X1 port map( A1 => n6687, A2 => n8860, B1 => n6879, B2 => 
                           n8857, ZN => n2612);
   U1667 : OAI22_X1 port map( A1 => n6688, A2 => n8860, B1 => n6880, B2 => 
                           n8857, ZN => n2630);
   U1668 : OAI22_X1 port map( A1 => n6689, A2 => n8860, B1 => n6881, B2 => 
                           n8857, ZN => n2648);
   U1669 : OAI22_X1 port map( A1 => n6690, A2 => n8860, B1 => n6882, B2 => 
                           n8857, ZN => n2666);
   U1670 : OAI22_X1 port map( A1 => n6691, A2 => n8859, B1 => n6883, B2 => 
                           n8856, ZN => n2684);
   U1671 : OAI22_X1 port map( A1 => n6692, A2 => n8859, B1 => n6884, B2 => 
                           n8856, ZN => n2702);
   U1672 : OAI22_X1 port map( A1 => n6693, A2 => n8859, B1 => n6885, B2 => 
                           n8856, ZN => n2720);
   U1673 : OAI22_X1 port map( A1 => n6694, A2 => n8859, B1 => n6886, B2 => 
                           n8856, ZN => n2738);
   U1674 : OAI22_X1 port map( A1 => n6695, A2 => n8859, B1 => n6887, B2 => 
                           n8856, ZN => n2756);
   U1675 : OAI22_X1 port map( A1 => n6696, A2 => n8859, B1 => n6888, B2 => 
                           n8856, ZN => n2774);
   U1676 : OAI22_X1 port map( A1 => n6697, A2 => n8859, B1 => n6889, B2 => 
                           n8856, ZN => n2792);
   U1677 : OAI22_X1 port map( A1 => n6698, A2 => n8859, B1 => n6890, B2 => 
                           n8856, ZN => n2810);
   U1678 : OAI22_X1 port map( A1 => n6699, A2 => n8859, B1 => n6891, B2 => 
                           n8856, ZN => n2828);
   U1679 : OAI22_X1 port map( A1 => n6700, A2 => n8859, B1 => n6892, B2 => 
                           n8856, ZN => n2846);
   U1680 : OAI22_X1 port map( A1 => n6701, A2 => n8859, B1 => n6893, B2 => 
                           n8856, ZN => n2864);
   U1681 : OAI22_X1 port map( A1 => n6702, A2 => n8859, B1 => n6894, B2 => 
                           n8856, ZN => n2882);
   U1682 : OAI22_X1 port map( A1 => n6703, A2 => n8858, B1 => n6895, B2 => 
                           n8855, ZN => n2900);
   U1683 : OAI22_X1 port map( A1 => n6704, A2 => n8858, B1 => n6896, B2 => 
                           n8855, ZN => n2918);
   U1684 : OAI22_X1 port map( A1 => n6705, A2 => n8858, B1 => n6897, B2 => 
                           n8855, ZN => n2936);
   U1685 : OAI22_X1 port map( A1 => n6706, A2 => n8858, B1 => n6898, B2 => 
                           n8855, ZN => n2954);
   U1686 : OAI22_X1 port map( A1 => n6667, A2 => n8858, B1 => n6859, B2 => 
                           n8855, ZN => n2972);
   U1687 : OAI22_X1 port map( A1 => n6668, A2 => n8858, B1 => n6860, B2 => 
                           n8855, ZN => n2990);
   U1688 : OAI22_X1 port map( A1 => n6669, A2 => n8858, B1 => n6861, B2 => 
                           n8855, ZN => n3008);
   U1689 : OAI22_X1 port map( A1 => n6670, A2 => n8858, B1 => n6862, B2 => 
                           n8855, ZN => n3026);
   U1690 : OAI22_X1 port map( A1 => n6671, A2 => n8858, B1 => n6863, B2 => 
                           n8855, ZN => n3044);
   U1691 : OAI22_X1 port map( A1 => n6672, A2 => n8858, B1 => n6864, B2 => 
                           n8855, ZN => n3062);
   U1692 : OAI22_X1 port map( A1 => n6673, A2 => n8858, B1 => n6865, B2 => 
                           n8855, ZN => n3080);
   U1693 : OAI22_X1 port map( A1 => n6674, A2 => n8858, B1 => n6866, B2 => 
                           n8855, ZN => n3109);
   U1694 : AOI22_X1 port map( A1 => n3815, A2 => n8989, B1 => n3671, B2 => 
                           n8986, ZN => n867);
   U1695 : AOI22_X1 port map( A1 => n3816, A2 => n8989, B1 => n3672, B2 => 
                           n8986, ZN => n908);
   U1696 : AOI22_X1 port map( A1 => n3817, A2 => n8989, B1 => n3673, B2 => 
                           n8986, ZN => n926);
   U1697 : AOI22_X1 port map( A1 => n3818, A2 => n8989, B1 => n3674, B2 => 
                           n8986, ZN => n944);
   U1698 : AOI22_X1 port map( A1 => n3819, A2 => n8989, B1 => n3675, B2 => 
                           n8986, ZN => n962);
   U1699 : AOI22_X1 port map( A1 => n3820, A2 => n8989, B1 => n3676, B2 => 
                           n8986, ZN => n980);
   U1700 : AOI22_X1 port map( A1 => n3821, A2 => n8989, B1 => n3677, B2 => 
                           n8986, ZN => n998);
   U1701 : AOI22_X1 port map( A1 => n3822, A2 => n8989, B1 => n3678, B2 => 
                           n8986, ZN => n1016);
   U1702 : OAI221_X1 port map( B1 => n8944, B2 => n7789, C1 => n8941, C2 => 
                           n7997, A => n892, ZN => n877);
   U1703 : AOI22_X1 port map( A1 => n3384, A2 => n8938, B1 => n3359, B2 => 
                           n8935, ZN => n892);
   U1704 : OAI221_X1 port map( B1 => n9019, B2 => n7877, C1 => n9016, C2 => 
                           n8157, A => n857, ZN => n854);
   U1705 : AOI22_X1 port map( A1 => n6635, A2 => n9013, B1 => n6347, B2 => 
                           n9010, ZN => n857);
   U1706 : OAI221_X1 port map( B1 => n8944, B2 => n7790, C1 => n8941, C2 => 
                           n7998, A => n916, ZN => n911);
   U1707 : AOI22_X1 port map( A1 => n3386, A2 => n8938, B1 => n3360, B2 => 
                           n8935, ZN => n916);
   U1708 : OAI221_X1 port map( B1 => n9019, B2 => n7878, C1 => n9016, C2 => 
                           n8158, A => n906, ZN => n905);
   U1709 : AOI22_X1 port map( A1 => n6636, A2 => n9013, B1 => n6348, B2 => 
                           n9010, ZN => n906);
   U1710 : OAI221_X1 port map( B1 => n8944, B2 => n7791, C1 => n8941, C2 => 
                           n7999, A => n934, ZN => n929);
   U1711 : AOI22_X1 port map( A1 => n3388, A2 => n8938, B1 => n3361, B2 => 
                           n8935, ZN => n934);
   U1712 : OAI221_X1 port map( B1 => n9019, B2 => n7879, C1 => n9016, C2 => 
                           n8159, A => n924, ZN => n923);
   U1713 : AOI22_X1 port map( A1 => n6637, A2 => n9013, B1 => n6349, B2 => 
                           n9010, ZN => n924);
   U1714 : OAI221_X1 port map( B1 => n8944, B2 => n7792, C1 => n8941, C2 => 
                           n8000, A => n952, ZN => n947);
   U1715 : AOI22_X1 port map( A1 => n3390, A2 => n8938, B1 => n3362, B2 => 
                           n8935, ZN => n952);
   U1716 : OAI221_X1 port map( B1 => n9019, B2 => n7880, C1 => n9016, C2 => 
                           n8160, A => n942, ZN => n941);
   U1717 : AOI22_X1 port map( A1 => n6638, A2 => n9013, B1 => n6350, B2 => 
                           n9010, ZN => n942);
   U1718 : OAI221_X1 port map( B1 => n8944, B2 => n7793, C1 => n8941, C2 => 
                           n8001, A => n970, ZN => n965);
   U1719 : AOI22_X1 port map( A1 => n3392, A2 => n8938, B1 => n3363, B2 => 
                           n8935, ZN => n970);
   U1720 : OAI221_X1 port map( B1 => n9019, B2 => n7881, C1 => n9016, C2 => 
                           n8161, A => n960, ZN => n959);
   U1721 : AOI22_X1 port map( A1 => n6639, A2 => n9013, B1 => n6351, B2 => 
                           n9010, ZN => n960);
   U1722 : OAI221_X1 port map( B1 => n8944, B2 => n7794, C1 => n8941, C2 => 
                           n8002, A => n988, ZN => n983);
   U1723 : AOI22_X1 port map( A1 => n3394, A2 => n8938, B1 => n3364, B2 => 
                           n8935, ZN => n988);
   U1724 : OAI221_X1 port map( B1 => n9019, B2 => n7882, C1 => n9016, C2 => 
                           n8162, A => n978, ZN => n977);
   U1725 : AOI22_X1 port map( A1 => n6640, A2 => n9013, B1 => n6352, B2 => 
                           n9010, ZN => n978);
   U1726 : OAI221_X1 port map( B1 => n8944, B2 => n7795, C1 => n8941, C2 => 
                           n8003, A => n1006, ZN => n1001);
   U1727 : AOI22_X1 port map( A1 => n3396, A2 => n8938, B1 => n3365, B2 => 
                           n8935, ZN => n1006);
   U1728 : OAI221_X1 port map( B1 => n9019, B2 => n7883, C1 => n9016, C2 => 
                           n8163, A => n996, ZN => n995);
   U1729 : AOI22_X1 port map( A1 => n6641, A2 => n9013, B1 => n6353, B2 => 
                           n9010, ZN => n996);
   U1730 : OAI221_X1 port map( B1 => n8944, B2 => n7796, C1 => n8941, C2 => 
                           n8004, A => n1024, ZN => n1019);
   U1731 : AOI22_X1 port map( A1 => n3398, A2 => n8938, B1 => n3366, B2 => 
                           n8935, ZN => n1024);
   U1732 : OAI221_X1 port map( B1 => n9019, B2 => n7884, C1 => n9016, C2 => 
                           n8164, A => n1014, ZN => n1013);
   U1733 : AOI22_X1 port map( A1 => n6642, A2 => n9013, B1 => n6354, B2 => 
                           n9010, ZN => n1014);
   U1734 : OAI22_X1 port map( A1 => n8452, A2 => n8791, B1 => n6619, B2 => 
                           n3189, ZN => n1328);
   U1735 : OAI22_X1 port map( A1 => n8453, A2 => n8794, B1 => n6620, B2 => 
                           n3189, ZN => n1329);
   U1736 : OAI22_X1 port map( A1 => n8453, A2 => n8797, B1 => n6621, B2 => 
                           n3189, ZN => n1330);
   U1737 : OAI22_X1 port map( A1 => n8453, A2 => n8800, B1 => n6622, B2 => 
                           n3189, ZN => n1331);
   U1738 : OAI22_X1 port map( A1 => n8453, A2 => n8803, B1 => n6623, B2 => 
                           n3189, ZN => n1332);
   U1739 : OAI22_X1 port map( A1 => n8453, A2 => n8806, B1 => n6624, B2 => 
                           n3189, ZN => n1333);
   U1740 : OAI22_X1 port map( A1 => n8454, A2 => n8809, B1 => n6625, B2 => 
                           n3189, ZN => n1334);
   U1741 : OAI22_X1 port map( A1 => n8454, A2 => n8821, B1 => n6626, B2 => 
                           n3189, ZN => n1335);
   U1742 : OAI22_X1 port map( A1 => n8461, A2 => n8791, B1 => n7941, B2 => 
                           n3188, ZN => n1360);
   U1743 : OAI22_X1 port map( A1 => n8462, A2 => n8794, B1 => n7942, B2 => 
                           n3188, ZN => n1361);
   U1744 : OAI22_X1 port map( A1 => n8462, A2 => n8797, B1 => n7943, B2 => 
                           n3188, ZN => n1362);
   U1745 : OAI22_X1 port map( A1 => n8462, A2 => n8800, B1 => n7944, B2 => 
                           n3188, ZN => n1363);
   U1746 : OAI22_X1 port map( A1 => n8462, A2 => n8803, B1 => n7945, B2 => 
                           n3188, ZN => n1364);
   U1747 : OAI22_X1 port map( A1 => n8462, A2 => n8806, B1 => n7946, B2 => 
                           n3188, ZN => n1365);
   U1748 : OAI22_X1 port map( A1 => n8463, A2 => n8809, B1 => n7947, B2 => 
                           n3188, ZN => n1366);
   U1749 : OAI22_X1 port map( A1 => n8463, A2 => n8821, B1 => n7948, B2 => 
                           n3188, ZN => n1367);
   U1750 : OAI22_X1 port map( A1 => n8470, A2 => n8791, B1 => n7949, B2 => 
                           n3187, ZN => n1392);
   U1751 : OAI22_X1 port map( A1 => n8471, A2 => n8794, B1 => n7950, B2 => 
                           n3187, ZN => n1393);
   U1752 : OAI22_X1 port map( A1 => n8471, A2 => n8797, B1 => n7951, B2 => 
                           n3187, ZN => n1394);
   U1753 : OAI22_X1 port map( A1 => n8471, A2 => n8800, B1 => n7952, B2 => 
                           n3187, ZN => n1395);
   U1754 : OAI22_X1 port map( A1 => n8471, A2 => n8803, B1 => n7953, B2 => 
                           n3187, ZN => n1396);
   U1755 : OAI22_X1 port map( A1 => n8471, A2 => n8806, B1 => n7954, B2 => 
                           n3187, ZN => n1397);
   U1756 : OAI22_X1 port map( A1 => n8472, A2 => n8809, B1 => n7955, B2 => 
                           n3187, ZN => n1398);
   U1757 : OAI22_X1 port map( A1 => n8472, A2 => n8821, B1 => n7956, B2 => 
                           n3187, ZN => n1399);
   U1758 : OAI22_X1 port map( A1 => n8488, A2 => n8791, B1 => n6667, B2 => 
                           n3185, ZN => n1456);
   U1759 : OAI22_X1 port map( A1 => n8489, A2 => n8794, B1 => n6668, B2 => 
                           n3185, ZN => n1457);
   U1760 : OAI22_X1 port map( A1 => n8489, A2 => n8797, B1 => n6669, B2 => 
                           n3185, ZN => n1458);
   U1761 : OAI22_X1 port map( A1 => n8489, A2 => n8800, B1 => n6670, B2 => 
                           n3185, ZN => n1459);
   U1762 : OAI22_X1 port map( A1 => n8489, A2 => n8803, B1 => n6671, B2 => 
                           n3185, ZN => n1460);
   U1763 : OAI22_X1 port map( A1 => n8489, A2 => n8806, B1 => n6672, B2 => 
                           n3185, ZN => n1461);
   U1764 : OAI22_X1 port map( A1 => n8490, A2 => n8809, B1 => n6673, B2 => 
                           n3185, ZN => n1462);
   U1765 : OAI22_X1 port map( A1 => n8490, A2 => n8821, B1 => n6674, B2 => 
                           n3185, ZN => n1463);
   U1766 : OAI22_X1 port map( A1 => n8506, A2 => n8791, B1 => n6859, B2 => 
                           n3182, ZN => n1520);
   U1767 : OAI22_X1 port map( A1 => n8507, A2 => n8794, B1 => n6860, B2 => 
                           n3182, ZN => n1521);
   U1768 : OAI22_X1 port map( A1 => n8507, A2 => n8797, B1 => n6861, B2 => 
                           n3182, ZN => n1522);
   U1769 : OAI22_X1 port map( A1 => n8507, A2 => n8800, B1 => n6862, B2 => 
                           n3182, ZN => n1523);
   U1770 : OAI22_X1 port map( A1 => n8507, A2 => n8803, B1 => n6863, B2 => 
                           n3182, ZN => n1524);
   U1771 : OAI22_X1 port map( A1 => n8507, A2 => n8806, B1 => n6864, B2 => 
                           n3182, ZN => n1525);
   U1772 : OAI22_X1 port map( A1 => n8508, A2 => n8809, B1 => n6865, B2 => 
                           n3182, ZN => n1526);
   U1773 : OAI22_X1 port map( A1 => n8508, A2 => n8821, B1 => n6866, B2 => 
                           n3182, ZN => n1527);
   U1774 : OAI22_X1 port map( A1 => n8515, A2 => n8790, B1 => n7925, B2 => 
                           n3181, ZN => n1552);
   U1775 : OAI22_X1 port map( A1 => n8516, A2 => n8793, B1 => n7926, B2 => 
                           n3181, ZN => n1553);
   U1776 : OAI22_X1 port map( A1 => n8516, A2 => n8796, B1 => n7927, B2 => 
                           n3181, ZN => n1554);
   U1777 : OAI22_X1 port map( A1 => n8516, A2 => n8799, B1 => n7928, B2 => 
                           n3181, ZN => n1555);
   U1778 : OAI22_X1 port map( A1 => n8516, A2 => n8802, B1 => n7929, B2 => 
                           n3181, ZN => n1556);
   U1779 : OAI22_X1 port map( A1 => n8516, A2 => n8805, B1 => n7930, B2 => 
                           n3181, ZN => n1557);
   U1780 : OAI22_X1 port map( A1 => n8517, A2 => n8808, B1 => n7931, B2 => 
                           n3181, ZN => n1558);
   U1781 : OAI22_X1 port map( A1 => n8517, A2 => n8820, B1 => n7932, B2 => 
                           n3181, ZN => n1559);
   U1782 : OAI22_X1 port map( A1 => n8533, A2 => n8790, B1 => n6331, B2 => 
                           n3179, ZN => n1616);
   U1783 : OAI22_X1 port map( A1 => n8534, A2 => n8793, B1 => n6332, B2 => 
                           n3179, ZN => n1617);
   U1784 : OAI22_X1 port map( A1 => n8534, A2 => n8796, B1 => n6333, B2 => 
                           n3179, ZN => n1618);
   U1785 : OAI22_X1 port map( A1 => n8534, A2 => n8799, B1 => n6334, B2 => 
                           n3179, ZN => n1619);
   U1786 : OAI22_X1 port map( A1 => n8534, A2 => n8802, B1 => n6335, B2 => 
                           n3179, ZN => n1620);
   U1787 : OAI22_X1 port map( A1 => n8534, A2 => n8805, B1 => n6336, B2 => 
                           n3179, ZN => n1621);
   U1788 : OAI22_X1 port map( A1 => n8535, A2 => n8808, B1 => n6337, B2 => 
                           n3179, ZN => n1622);
   U1789 : OAI22_X1 port map( A1 => n8535, A2 => n8820, B1 => n6338, B2 => 
                           n3179, ZN => n1623);
   U1790 : OAI22_X1 port map( A1 => n8551, A2 => n8790, B1 => n7933, B2 => 
                           n3177, ZN => n1680);
   U1791 : OAI22_X1 port map( A1 => n8552, A2 => n8793, B1 => n7934, B2 => 
                           n3177, ZN => n1681);
   U1792 : OAI22_X1 port map( A1 => n8552, A2 => n8796, B1 => n7935, B2 => 
                           n3177, ZN => n1682);
   U1793 : OAI22_X1 port map( A1 => n8552, A2 => n8799, B1 => n7936, B2 => 
                           n3177, ZN => n1683);
   U1794 : OAI22_X1 port map( A1 => n8552, A2 => n8802, B1 => n7937, B2 => 
                           n3177, ZN => n1684);
   U1795 : OAI22_X1 port map( A1 => n8552, A2 => n8805, B1 => n7938, B2 => 
                           n3177, ZN => n1685);
   U1796 : OAI22_X1 port map( A1 => n8553, A2 => n8808, B1 => n7939, B2 => 
                           n3177, ZN => n1686);
   U1797 : OAI22_X1 port map( A1 => n8553, A2 => n8820, B1 => n7940, B2 => 
                           n3177, ZN => n1687);
   U1798 : OAI22_X1 port map( A1 => n8560, A2 => n8790, B1 => n6675, B2 => 
                           n3176, ZN => n1712);
   U1799 : OAI22_X1 port map( A1 => n8561, A2 => n8793, B1 => n6676, B2 => 
                           n3176, ZN => n1713);
   U1800 : OAI22_X1 port map( A1 => n8561, A2 => n8796, B1 => n6677, B2 => 
                           n3176, ZN => n1714);
   U1801 : OAI22_X1 port map( A1 => n8561, A2 => n8799, B1 => n6678, B2 => 
                           n3176, ZN => n1715);
   U1802 : OAI22_X1 port map( A1 => n8561, A2 => n8802, B1 => n6679, B2 => 
                           n3176, ZN => n1716);
   U1803 : OAI22_X1 port map( A1 => n8561, A2 => n8805, B1 => n6680, B2 => 
                           n3176, ZN => n1717);
   U1804 : OAI22_X1 port map( A1 => n8562, A2 => n8808, B1 => n6681, B2 => 
                           n3176, ZN => n1718);
   U1805 : OAI22_X1 port map( A1 => n8562, A2 => n8820, B1 => n6682, B2 => 
                           n3176, ZN => n1719);
   U1806 : OAI22_X1 port map( A1 => n8596, A2 => n8790, B1 => n6795, B2 => 
                           n3171, ZN => n1840);
   U1807 : OAI22_X1 port map( A1 => n8597, A2 => n8793, B1 => n6796, B2 => 
                           n3171, ZN => n1841);
   U1808 : OAI22_X1 port map( A1 => n8597, A2 => n8796, B1 => n6797, B2 => 
                           n3171, ZN => n1842);
   U1809 : OAI22_X1 port map( A1 => n8597, A2 => n8799, B1 => n6798, B2 => 
                           n3171, ZN => n1843);
   U1810 : OAI22_X1 port map( A1 => n8597, A2 => n8802, B1 => n6799, B2 => 
                           n3171, ZN => n1844);
   U1811 : OAI22_X1 port map( A1 => n8597, A2 => n8805, B1 => n6800, B2 => 
                           n3171, ZN => n1845);
   U1812 : OAI22_X1 port map( A1 => n8598, A2 => n8808, B1 => n6801, B2 => 
                           n3171, ZN => n1846);
   U1813 : OAI22_X1 port map( A1 => n8598, A2 => n8820, B1 => n6802, B2 => 
                           n3171, ZN => n1847);
   U1814 : OAI22_X1 port map( A1 => n8605, A2 => n8790, B1 => n6731, B2 => 
                           n3170, ZN => n1872);
   U1815 : OAI22_X1 port map( A1 => n8606, A2 => n8793, B1 => n6732, B2 => 
                           n3170, ZN => n1873);
   U1816 : OAI22_X1 port map( A1 => n8606, A2 => n8796, B1 => n6733, B2 => 
                           n3170, ZN => n1874);
   U1817 : OAI22_X1 port map( A1 => n8606, A2 => n8799, B1 => n6734, B2 => 
                           n3170, ZN => n1875);
   U1818 : OAI22_X1 port map( A1 => n8606, A2 => n8802, B1 => n6735, B2 => 
                           n3170, ZN => n1876);
   U1819 : OAI22_X1 port map( A1 => n8606, A2 => n8805, B1 => n6736, B2 => 
                           n3170, ZN => n1877);
   U1820 : OAI22_X1 port map( A1 => n8607, A2 => n8808, B1 => n6737, B2 => 
                           n3170, ZN => n1878);
   U1821 : OAI22_X1 port map( A1 => n8607, A2 => n8820, B1 => n6738, B2 => 
                           n3170, ZN => n1879);
   U1822 : OAI22_X1 port map( A1 => n8614, A2 => n8790, B1 => n6739, B2 => 
                           n3169, ZN => n1904);
   U1823 : OAI22_X1 port map( A1 => n8615, A2 => n8793, B1 => n6740, B2 => 
                           n3169, ZN => n1905);
   U1824 : OAI22_X1 port map( A1 => n8615, A2 => n8796, B1 => n6741, B2 => 
                           n3169, ZN => n1906);
   U1825 : OAI22_X1 port map( A1 => n8615, A2 => n8799, B1 => n6742, B2 => 
                           n3169, ZN => n1907);
   U1826 : OAI22_X1 port map( A1 => n8615, A2 => n8802, B1 => n6743, B2 => 
                           n3169, ZN => n1908);
   U1827 : OAI22_X1 port map( A1 => n8615, A2 => n8805, B1 => n6744, B2 => 
                           n3169, ZN => n1909);
   U1828 : OAI22_X1 port map( A1 => n8616, A2 => n8808, B1 => n6745, B2 => 
                           n3169, ZN => n1910);
   U1829 : OAI22_X1 port map( A1 => n8616, A2 => n8820, B1 => n6746, B2 => 
                           n3169, ZN => n1911);
   U1830 : OAI22_X1 port map( A1 => n8623, A2 => n8789, B1 => n7957, B2 => 
                           n3168, ZN => n1936);
   U1831 : OAI22_X1 port map( A1 => n8624, A2 => n8792, B1 => n7958, B2 => 
                           n3168, ZN => n1937);
   U1832 : OAI22_X1 port map( A1 => n8624, A2 => n8795, B1 => n7959, B2 => 
                           n3168, ZN => n1938);
   U1833 : OAI22_X1 port map( A1 => n8624, A2 => n8798, B1 => n7960, B2 => 
                           n3168, ZN => n1939);
   U1834 : OAI22_X1 port map( A1 => n8624, A2 => n8801, B1 => n7961, B2 => 
                           n3168, ZN => n1940);
   U1835 : OAI22_X1 port map( A1 => n8624, A2 => n8804, B1 => n7962, B2 => 
                           n3168, ZN => n1941);
   U1836 : OAI22_X1 port map( A1 => n8625, A2 => n8807, B1 => n7963, B2 => 
                           n3168, ZN => n1942);
   U1837 : OAI22_X1 port map( A1 => n8625, A2 => n8819, B1 => n7964, B2 => 
                           n3168, ZN => n1943);
   U1838 : OAI22_X1 port map( A1 => n8641, A2 => n8789, B1 => n6867, B2 => 
                           n3166, ZN => n2000);
   U1839 : OAI22_X1 port map( A1 => n8642, A2 => n8792, B1 => n6868, B2 => 
                           n3166, ZN => n2001);
   U1840 : OAI22_X1 port map( A1 => n8642, A2 => n8795, B1 => n6869, B2 => 
                           n3166, ZN => n2002);
   U1841 : OAI22_X1 port map( A1 => n8642, A2 => n8798, B1 => n6870, B2 => 
                           n3166, ZN => n2003);
   U1842 : OAI22_X1 port map( A1 => n8642, A2 => n8801, B1 => n6871, B2 => 
                           n3166, ZN => n2004);
   U1843 : OAI22_X1 port map( A1 => n8642, A2 => n8804, B1 => n6872, B2 => 
                           n3166, ZN => n2005);
   U1844 : OAI22_X1 port map( A1 => n8643, A2 => n8807, B1 => n6873, B2 => 
                           n3166, ZN => n2006);
   U1845 : OAI22_X1 port map( A1 => n8643, A2 => n8819, B1 => n6874, B2 => 
                           n3166, ZN => n2007);
   U1846 : OAI22_X1 port map( A1 => n8677, A2 => n8789, B1 => n6803, B2 => 
                           n3158, ZN => n2128);
   U1847 : OAI22_X1 port map( A1 => n8678, A2 => n8792, B1 => n6804, B2 => 
                           n3158, ZN => n2129);
   U1848 : OAI22_X1 port map( A1 => n8678, A2 => n8795, B1 => n6805, B2 => 
                           n3158, ZN => n2130);
   U1849 : OAI22_X1 port map( A1 => n8678, A2 => n8798, B1 => n6806, B2 => 
                           n3158, ZN => n2131);
   U1850 : OAI22_X1 port map( A1 => n8678, A2 => n8801, B1 => n6807, B2 => 
                           n3158, ZN => n2132);
   U1851 : OAI22_X1 port map( A1 => n8678, A2 => n8804, B1 => n6808, B2 => 
                           n3158, ZN => n2133);
   U1852 : OAI22_X1 port map( A1 => n8679, A2 => n8807, B1 => n6809, B2 => 
                           n3158, ZN => n2134);
   U1853 : OAI22_X1 port map( A1 => n8679, A2 => n8819, B1 => n6810, B2 => 
                           n3158, ZN => n2135);
   U1854 : OAI22_X1 port map( A1 => n8686, A2 => n8789, B1 => n7965, B2 => 
                           n3156, ZN => n2160);
   U1855 : OAI22_X1 port map( A1 => n8687, A2 => n8792, B1 => n7966, B2 => 
                           n3156, ZN => n2161);
   U1856 : OAI22_X1 port map( A1 => n8687, A2 => n8795, B1 => n7967, B2 => 
                           n3156, ZN => n2162);
   U1857 : OAI22_X1 port map( A1 => n8687, A2 => n8798, B1 => n7968, B2 => 
                           n3156, ZN => n2163);
   U1858 : OAI22_X1 port map( A1 => n8687, A2 => n8801, B1 => n7969, B2 => 
                           n3156, ZN => n2164);
   U1859 : OAI22_X1 port map( A1 => n8687, A2 => n8804, B1 => n7970, B2 => 
                           n3156, ZN => n2165);
   U1860 : OAI22_X1 port map( A1 => n8688, A2 => n8807, B1 => n7971, B2 => 
                           n3156, ZN => n2166);
   U1861 : OAI22_X1 port map( A1 => n8688, A2 => n8819, B1 => n7972, B2 => 
                           n3156, ZN => n2167);
   U1862 : AOI22_X1 port map( A1 => n3823, A2 => n8988, B1 => n3679, B2 => 
                           n8985, ZN => n1034);
   U1863 : AOI22_X1 port map( A1 => n3824, A2 => n8988, B1 => n3680, B2 => 
                           n8985, ZN => n1052);
   U1864 : AOI22_X1 port map( A1 => n3825, A2 => n8988, B1 => n3681, B2 => 
                           n8985, ZN => n1070);
   U1865 : AOI22_X1 port map( A1 => n3826, A2 => n8988, B1 => n3682, B2 => 
                           n8985, ZN => n1088);
   U1866 : AOI22_X1 port map( A1 => n3827, A2 => n8988, B1 => n3683, B2 => 
                           n8985, ZN => n1106);
   U1867 : AOI22_X1 port map( A1 => n3828, A2 => n8988, B1 => n3684, B2 => 
                           n8985, ZN => n1124);
   U1868 : AOI22_X1 port map( A1 => n3829, A2 => n8988, B1 => n3685, B2 => 
                           n8985, ZN => n1142);
   U1869 : AOI22_X1 port map( A1 => n3830, A2 => n8988, B1 => n3686, B2 => 
                           n8985, ZN => n1160);
   U1870 : AOI22_X1 port map( A1 => n3831, A2 => n8988, B1 => n3687, B2 => 
                           n8985, ZN => n1178);
   U1871 : AOI22_X1 port map( A1 => n3832, A2 => n8988, B1 => n3688, B2 => 
                           n8985, ZN => n1196);
   U1872 : AOI22_X1 port map( A1 => n3833, A2 => n8988, B1 => n3689, B2 => 
                           n8985, ZN => n1214);
   U1873 : AOI22_X1 port map( A1 => n3834, A2 => n8988, B1 => n3690, B2 => 
                           n8985, ZN => n1232);
   U1874 : AOI22_X1 port map( A1 => n3835, A2 => n8987, B1 => n3691, B2 => 
                           n8984, ZN => n1250);
   U1875 : AOI22_X1 port map( A1 => n3836, A2 => n8987, B1 => n3692, B2 => 
                           n8984, ZN => n1268);
   U1876 : AOI22_X1 port map( A1 => n3837, A2 => n8987, B1 => n3693, B2 => 
                           n8984, ZN => n2310);
   U1877 : AOI22_X1 port map( A1 => n3838, A2 => n8987, B1 => n3694, B2 => 
                           n8984, ZN => n2328);
   U1878 : AOI22_X1 port map( A1 => n3607, A2 => n8987, B1 => n3583, B2 => 
                           n8984, ZN => n2346);
   U1879 : AOI22_X1 port map( A1 => n3608, A2 => n8987, B1 => n3584, B2 => 
                           n8984, ZN => n2364);
   U1880 : AOI22_X1 port map( A1 => n3609, A2 => n8987, B1 => n3585, B2 => 
                           n8984, ZN => n2382);
   U1881 : AOI22_X1 port map( A1 => n3610, A2 => n8987, B1 => n3586, B2 => 
                           n8984, ZN => n2400);
   U1882 : AOI22_X1 port map( A1 => n3611, A2 => n8987, B1 => n3587, B2 => 
                           n8984, ZN => n2418);
   U1883 : AOI22_X1 port map( A1 => n3612, A2 => n8987, B1 => n3588, B2 => 
                           n8984, ZN => n2436);
   U1884 : AOI22_X1 port map( A1 => n3613, A2 => n8987, B1 => n3589, B2 => 
                           n8984, ZN => n2454);
   U1885 : AOI22_X1 port map( A1 => n3614, A2 => n8987, B1 => n3590, B2 => 
                           n8984, ZN => n2481);
   U1886 : AOI22_X1 port map( A1 => n8914, A2 => n8053, B1 => n8910, B2 => 
                           OUT1_0_port, ZN => n2504);
   U1887 : AOI22_X1 port map( A1 => n8890, A2 => n3384, B1 => n8885, B2 => 
                           n3359, ZN => n2514);
   U1888 : AOI22_X1 port map( A1 => n8878, A2 => n3479, B1 => n8873, B2 => 
                           n3767, ZN => n2519);
   U1889 : AOI22_X1 port map( A1 => n8914, A2 => n8054, B1 => n8909, B2 => 
                           OUT1_1_port, ZN => n2553);
   U1890 : AOI22_X1 port map( A1 => n8890, A2 => n3386, B1 => n8885, B2 => 
                           n3360, ZN => n2555);
   U1891 : AOI22_X1 port map( A1 => n8878, A2 => n3480, B1 => n8873, B2 => 
                           n3768, ZN => n2556);
   U1892 : AOI22_X1 port map( A1 => n8914, A2 => n8055, B1 => n8909, B2 => 
                           OUT1_2_port, ZN => n2571);
   U1893 : AOI22_X1 port map( A1 => n8890, A2 => n3388, B1 => n8885, B2 => 
                           n3361, ZN => n2573);
   U1894 : AOI22_X1 port map( A1 => n8878, A2 => n3481, B1 => n8873, B2 => 
                           n3769, ZN => n2574);
   U1895 : AOI22_X1 port map( A1 => n8914, A2 => n8056, B1 => n8909, B2 => 
                           OUT1_3_port, ZN => n2589);
   U1896 : AOI22_X1 port map( A1 => n8890, A2 => n3390, B1 => n8885, B2 => 
                           n3362, ZN => n2591);
   U1897 : AOI22_X1 port map( A1 => n8878, A2 => n3482, B1 => n8873, B2 => 
                           n3770, ZN => n2592);
   U1898 : AOI22_X1 port map( A1 => n8914, A2 => n8057, B1 => n8909, B2 => 
                           OUT1_4_port, ZN => n2607);
   U1899 : AOI22_X1 port map( A1 => n8890, A2 => n3392, B1 => n8885, B2 => 
                           n3363, ZN => n2609);
   U1900 : AOI22_X1 port map( A1 => n8878, A2 => n3483, B1 => n8873, B2 => 
                           n3771, ZN => n2610);
   U1901 : AOI22_X1 port map( A1 => n8914, A2 => n8058, B1 => n8909, B2 => 
                           OUT1_5_port, ZN => n2625);
   U1902 : AOI22_X1 port map( A1 => n8890, A2 => n3394, B1 => n8885, B2 => 
                           n3364, ZN => n2627);
   U1903 : AOI22_X1 port map( A1 => n8878, A2 => n3484, B1 => n8873, B2 => 
                           n3772, ZN => n2628);
   U1904 : AOI22_X1 port map( A1 => n8914, A2 => n8059, B1 => n8909, B2 => 
                           OUT1_6_port, ZN => n2643);
   U1905 : AOI22_X1 port map( A1 => n8890, A2 => n3396, B1 => n8885, B2 => 
                           n3365, ZN => n2645);
   U1906 : AOI22_X1 port map( A1 => n8878, A2 => n3485, B1 => n8873, B2 => 
                           n3773, ZN => n2646);
   U1907 : AOI22_X1 port map( A1 => n8914, A2 => n8060, B1 => n8909, B2 => 
                           OUT1_7_port, ZN => n2661);
   U1908 : AOI22_X1 port map( A1 => n8890, A2 => n3398, B1 => n8885, B2 => 
                           n3366, ZN => n2663);
   U1909 : AOI22_X1 port map( A1 => n8878, A2 => n3486, B1 => n8873, B2 => 
                           n3774, ZN => n2664);
   U1910 : AOI22_X1 port map( A1 => n8913, A2 => n8061, B1 => n8909, B2 => 
                           OUT1_8_port, ZN => n2679);
   U1911 : AOI22_X1 port map( A1 => n8889, A2 => n3400, B1 => n8885, B2 => 
                           n3367, ZN => n2681);
   U1912 : AOI22_X1 port map( A1 => n8877, A2 => n3519, B1 => n8873, B2 => 
                           n3775, ZN => n2682);
   U1913 : AOI22_X1 port map( A1 => n8913, A2 => n8062, B1 => n8910, B2 => 
                           OUT1_9_port, ZN => n2697);
   U1914 : AOI22_X1 port map( A1 => n8889, A2 => n3402, B1 => n8885, B2 => 
                           n3368, ZN => n2699);
   U1915 : AOI22_X1 port map( A1 => n8877, A2 => n3520, B1 => n8873, B2 => 
                           n3776, ZN => n2700);
   U1916 : AOI22_X1 port map( A1 => n8913, A2 => n8063, B1 => n8910, B2 => 
                           OUT1_10_port, ZN => n2715);
   U1917 : AOI22_X1 port map( A1 => n8889, A2 => n3404, B1 => n8885, B2 => 
                           n3369, ZN => n2717);
   U1918 : AOI22_X1 port map( A1 => n8877, A2 => n3521, B1 => n8873, B2 => 
                           n3777, ZN => n2718);
   U1919 : AOI22_X1 port map( A1 => n8913, A2 => n8064, B1 => n8910, B2 => 
                           OUT1_11_port, ZN => n2733);
   U1920 : AOI22_X1 port map( A1 => n8889, A2 => n3406, B1 => n8885, B2 => 
                           n3370, ZN => n2735);
   U1921 : AOI22_X1 port map( A1 => n8877, A2 => n3522, B1 => n8873, B2 => 
                           n3778, ZN => n2736);
   U1922 : AOI22_X1 port map( A1 => n8913, A2 => n8065, B1 => n8910, B2 => 
                           OUT1_12_port, ZN => n2751);
   U1923 : AOI22_X1 port map( A1 => n8889, A2 => n3408, B1 => n8886, B2 => 
                           n3371, ZN => n2753);
   U1924 : AOI22_X1 port map( A1 => n8877, A2 => n3523, B1 => n8874, B2 => 
                           n3779, ZN => n2754);
   U1925 : AOI22_X1 port map( A1 => n8913, A2 => n8066, B1 => n8910, B2 => 
                           OUT1_13_port, ZN => n2769);
   U1926 : AOI22_X1 port map( A1 => n8889, A2 => n3410, B1 => n8886, B2 => 
                           n3372, ZN => n2771);
   U1927 : AOI22_X1 port map( A1 => n8877, A2 => n3524, B1 => n8874, B2 => 
                           n3780, ZN => n2772);
   U1928 : AOI22_X1 port map( A1 => n8913, A2 => n8067, B1 => n8910, B2 => 
                           OUT1_14_port, ZN => n2787);
   U1929 : AOI22_X1 port map( A1 => n8889, A2 => n3412, B1 => n8886, B2 => 
                           n3373, ZN => n2789);
   U1930 : AOI22_X1 port map( A1 => n8877, A2 => n3525, B1 => n8874, B2 => 
                           n3781, ZN => n2790);
   U1931 : AOI22_X1 port map( A1 => n8913, A2 => n8068, B1 => n8910, B2 => 
                           OUT1_15_port, ZN => n2805);
   U1932 : AOI22_X1 port map( A1 => n8889, A2 => n3414, B1 => n8886, B2 => 
                           n3374, ZN => n2807);
   U1933 : AOI22_X1 port map( A1 => n8877, A2 => n3526, B1 => n8874, B2 => 
                           n3782, ZN => n2808);
   U1934 : AOI22_X1 port map( A1 => n8913, A2 => n8069, B1 => n8910, B2 => 
                           OUT1_16_port, ZN => n2823);
   U1935 : AOI22_X1 port map( A1 => n8889, A2 => n3416, B1 => n8886, B2 => 
                           n3375, ZN => n2825);
   U1936 : AOI22_X1 port map( A1 => n8877, A2 => n3527, B1 => n8874, B2 => 
                           n3783, ZN => n2826);
   U1937 : AOI22_X1 port map( A1 => n8913, A2 => n8070, B1 => n8910, B2 => 
                           OUT1_17_port, ZN => n2841);
   U1938 : AOI22_X1 port map( A1 => n8889, A2 => n3418, B1 => n8886, B2 => 
                           n3376, ZN => n2843);
   U1939 : AOI22_X1 port map( A1 => n8877, A2 => n3528, B1 => n8874, B2 => 
                           n3784, ZN => n2844);
   U1940 : AOI22_X1 port map( A1 => n8913, A2 => n8071, B1 => n8910, B2 => 
                           OUT1_18_port, ZN => n2859);
   U1941 : AOI22_X1 port map( A1 => n8889, A2 => n3420, B1 => n8886, B2 => 
                           n3377, ZN => n2861);
   U1942 : AOI22_X1 port map( A1 => n8877, A2 => n3529, B1 => n8874, B2 => 
                           n3785, ZN => n2862);
   U1943 : AOI22_X1 port map( A1 => n8913, A2 => n8072, B1 => n8910, B2 => 
                           OUT1_19_port, ZN => n2877);
   U1944 : AOI22_X1 port map( A1 => n8889, A2 => n3422, B1 => n8886, B2 => 
                           n3378, ZN => n2879);
   U1945 : AOI22_X1 port map( A1 => n8877, A2 => n3530, B1 => n8874, B2 => 
                           n3786, ZN => n2880);
   U1946 : AOI22_X1 port map( A1 => n8912, A2 => n8073, B1 => n8910, B2 => 
                           OUT1_20_port, ZN => n2895);
   U1947 : AOI22_X1 port map( A1 => n8888, A2 => n3424, B1 => n8886, B2 => 
                           n3379, ZN => n2897);
   U1948 : AOI22_X1 port map( A1 => n8876, A2 => n3531, B1 => n8874, B2 => 
                           n3787, ZN => n2898);
   U1949 : AOI22_X1 port map( A1 => n8912, A2 => n8074, B1 => n8911, B2 => 
                           OUT1_21_port, ZN => n2913);
   U1950 : AOI22_X1 port map( A1 => n8888, A2 => n3426, B1 => n8886, B2 => 
                           n3380, ZN => n2915);
   U1951 : AOI22_X1 port map( A1 => n8876, A2 => n3532, B1 => n8874, B2 => 
                           n3788, ZN => n2916);
   U1952 : AOI22_X1 port map( A1 => n8912, A2 => n8075, B1 => n8911, B2 => 
                           OUT1_22_port, ZN => n2931);
   U1953 : AOI22_X1 port map( A1 => n8888, A2 => n3428, B1 => n8886, B2 => 
                           n3381, ZN => n2933);
   U1954 : AOI22_X1 port map( A1 => n8876, A2 => n3533, B1 => n8874, B2 => 
                           n3789, ZN => n2934);
   U1955 : AOI22_X1 port map( A1 => n8912, A2 => n8076, B1 => n8911, B2 => 
                           OUT1_23_port, ZN => n2949);
   U1956 : AOI22_X1 port map( A1 => n8888, A2 => n3430, B1 => n8886, B2 => 
                           n3382, ZN => n2951);
   U1957 : AOI22_X1 port map( A1 => n8876, A2 => n3534, B1 => n8874, B2 => 
                           n3790, ZN => n2952);
   U1958 : AOI22_X1 port map( A1 => n8912, A2 => n8077, B1 => n8911, B2 => 
                           OUT1_24_port, ZN => n2967);
   U1959 : AOI22_X1 port map( A1 => n8888, A2 => n3432, B1 => n8887, B2 => 
                           n3279, ZN => n2969);
   U1960 : AOI22_X1 port map( A1 => n8876, A2 => n3535, B1 => n8875, B2 => 
                           n3567, ZN => n2970);
   U1961 : AOI22_X1 port map( A1 => n8912, A2 => n8078, B1 => n8911, B2 => 
                           OUT1_25_port, ZN => n2985);
   U1962 : AOI22_X1 port map( A1 => n8888, A2 => n3434, B1 => n8887, B2 => 
                           n3280, ZN => n2987);
   U1963 : AOI22_X1 port map( A1 => n8876, A2 => n3536, B1 => n8875, B2 => 
                           n3568, ZN => n2988);
   U1964 : AOI22_X1 port map( A1 => n8912, A2 => n8079, B1 => n8911, B2 => 
                           OUT1_26_port, ZN => n3003);
   U1965 : AOI22_X1 port map( A1 => n8888, A2 => n3436, B1 => n8887, B2 => 
                           n3281, ZN => n3005);
   U1966 : AOI22_X1 port map( A1 => n8876, A2 => n3537, B1 => n8875, B2 => 
                           n3569, ZN => n3006);
   U1967 : AOI22_X1 port map( A1 => n8912, A2 => n8080, B1 => n8911, B2 => 
                           OUT1_27_port, ZN => n3021);
   U1968 : AOI22_X1 port map( A1 => n8888, A2 => n3438, B1 => n8887, B2 => 
                           n3282, ZN => n3023);
   U1969 : AOI22_X1 port map( A1 => n8876, A2 => n3538, B1 => n8875, B2 => 
                           n3570, ZN => n3024);
   U1970 : AOI22_X1 port map( A1 => n8912, A2 => n8081, B1 => n8911, B2 => 
                           OUT1_28_port, ZN => n3039);
   U1971 : AOI22_X1 port map( A1 => n8888, A2 => n3440, B1 => n8887, B2 => 
                           n3283, ZN => n3041);
   U1972 : AOI22_X1 port map( A1 => n8876, A2 => n3539, B1 => n8875, B2 => 
                           n3571, ZN => n3042);
   U1973 : AOI22_X1 port map( A1 => n8912, A2 => n8082, B1 => n8911, B2 => 
                           OUT1_29_port, ZN => n3057);
   U1974 : AOI22_X1 port map( A1 => n8888, A2 => n3442, B1 => n8887, B2 => 
                           n3284, ZN => n3059);
   U1975 : AOI22_X1 port map( A1 => n8876, A2 => n3540, B1 => n8875, B2 => 
                           n3572, ZN => n3060);
   U1976 : AOI22_X1 port map( A1 => n8912, A2 => n8083, B1 => n8911, B2 => 
                           OUT1_30_port, ZN => n3075);
   U1977 : AOI22_X1 port map( A1 => n8888, A2 => n3444, B1 => n8887, B2 => 
                           n3285, ZN => n3077);
   U1978 : AOI22_X1 port map( A1 => n8876, A2 => n3541, B1 => n8875, B2 => 
                           n3573, ZN => n3078);
   U1979 : AOI22_X1 port map( A1 => n8912, A2 => n8084, B1 => n8909, B2 => 
                           OUT1_31_port, ZN => n3093);
   U1980 : AOI22_X1 port map( A1 => n8888, A2 => n3446, B1 => n8887, B2 => 
                           n3286, ZN => n3101);
   U1981 : AOI22_X1 port map( A1 => n8876, A2 => n3542, B1 => n8875, B2 => 
                           n3574, ZN => n3104);
   U1982 : OAI221_X1 port map( B1 => n8968, B2 => n7973, C1 => n6747, C2 => 
                           n8965, A => n882, ZN => n879);
   U1983 : AOI22_X1 port map( A1 => n8962, A2 => n8053, B1 => n8958, B2 => 
                           OUT2_0_port, ZN => n882);
   U1984 : OAI221_X1 port map( B1 => n8968, B2 => n7974, C1 => n6748, C2 => 
                           n8965, A => n914, ZN => n913);
   U1985 : AOI22_X1 port map( A1 => n8962, A2 => n8054, B1 => n8957, B2 => 
                           OUT2_1_port, ZN => n914);
   U1986 : OAI221_X1 port map( B1 => n8968, B2 => n7975, C1 => n6749, C2 => 
                           n8965, A => n932, ZN => n931);
   U1987 : AOI22_X1 port map( A1 => n8962, A2 => n8055, B1 => n8957, B2 => 
                           OUT2_2_port, ZN => n932);
   U1988 : OAI221_X1 port map( B1 => n8968, B2 => n7976, C1 => n6750, C2 => 
                           n8965, A => n950, ZN => n949);
   U1989 : AOI22_X1 port map( A1 => n8962, A2 => n8056, B1 => n8957, B2 => 
                           OUT2_3_port, ZN => n950);
   U1990 : OAI221_X1 port map( B1 => n8968, B2 => n7977, C1 => n6751, C2 => 
                           n8965, A => n968, ZN => n967);
   U1991 : AOI22_X1 port map( A1 => n8962, A2 => n8057, B1 => n8957, B2 => 
                           OUT2_4_port, ZN => n968);
   U1992 : OAI221_X1 port map( B1 => n8968, B2 => n7978, C1 => n6752, C2 => 
                           n8965, A => n986, ZN => n985);
   U1993 : AOI22_X1 port map( A1 => n8962, A2 => n8058, B1 => n8957, B2 => 
                           OUT2_5_port, ZN => n986);
   U1994 : OAI221_X1 port map( B1 => n8968, B2 => n7979, C1 => n6753, C2 => 
                           n8965, A => n1004, ZN => n1003);
   U1995 : AOI22_X1 port map( A1 => n8962, A2 => n8059, B1 => n8957, B2 => 
                           OUT2_6_port, ZN => n1004);
   U1996 : OAI221_X1 port map( B1 => n8968, B2 => n7980, C1 => n6754, C2 => 
                           n8965, A => n1022, ZN => n1021);
   U1997 : AOI22_X1 port map( A1 => n8962, A2 => n8060, B1 => n8957, B2 => 
                           OUT2_7_port, ZN => n1022);
   U1998 : OAI221_X1 port map( B1 => n8955, B2 => n8141, C1 => n6779, C2 => 
                           n8952, A => n1041, ZN => n1038);
   U1999 : AOI22_X1 port map( A1 => n8949, A2 => n8237, B1 => n3319, B2 => 
                           n8946, ZN => n1041);
   U2000 : OAI221_X1 port map( B1 => n8967, B2 => n7981, C1 => n6755, C2 => 
                           n8964, A => n1040, ZN => n1039);
   U2001 : AOI22_X1 port map( A1 => n8961, A2 => n8061, B1 => n8957, B2 => 
                           OUT2_8_port, ZN => n1040);
   U2002 : OAI221_X1 port map( B1 => n8943, B2 => n7797, C1 => n8940, C2 => 
                           n8005, A => n1042, ZN => n1037);
   U2003 : AOI22_X1 port map( A1 => n3400, A2 => n8937, B1 => n3367, B2 => 
                           n8934, ZN => n1042);
   U2004 : OAI221_X1 port map( B1 => n8931, B2 => n7798, C1 => n8928, C2 => 
                           n8037, A => n1043, ZN => n1036);
   U2005 : AOI22_X1 port map( A1 => n3519, A2 => n8925, B1 => n3775, B2 => 
                           n8922, ZN => n1043);
   U2006 : OAI221_X1 port map( B1 => n9018, B2 => n7885, C1 => n9015, C2 => 
                           n8165, A => n1032, ZN => n1031);
   U2007 : AOI22_X1 port map( A1 => n6643, A2 => n9012, B1 => n6355, B2 => 
                           n9009, ZN => n1032);
   U2008 : OAI221_X1 port map( B1 => n8955, B2 => n8142, C1 => n6780, C2 => 
                           n8952, A => n1059, ZN => n1056);
   U2009 : AOI22_X1 port map( A1 => n8949, A2 => n8238, B1 => n3320, B2 => 
                           n8946, ZN => n1059);
   U2010 : OAI221_X1 port map( B1 => n8967, B2 => n7982, C1 => n6756, C2 => 
                           n8964, A => n1058, ZN => n1057);
   U2011 : AOI22_X1 port map( A1 => n8961, A2 => n8062, B1 => n8958, B2 => 
                           OUT2_9_port, ZN => n1058);
   U2012 : OAI221_X1 port map( B1 => n8943, B2 => n7799, C1 => n8940, C2 => 
                           n8006, A => n1060, ZN => n1055);
   U2013 : AOI22_X1 port map( A1 => n3402, A2 => n8937, B1 => n3368, B2 => 
                           n8934, ZN => n1060);
   U2014 : OAI221_X1 port map( B1 => n8931, B2 => n7800, C1 => n8928, C2 => 
                           n8038, A => n1061, ZN => n1054);
   U2015 : AOI22_X1 port map( A1 => n3520, A2 => n8925, B1 => n3776, B2 => 
                           n8922, ZN => n1061);
   U2016 : OAI221_X1 port map( B1 => n9018, B2 => n7886, C1 => n9015, C2 => 
                           n8166, A => n1050, ZN => n1049);
   U2017 : AOI22_X1 port map( A1 => n6644, A2 => n9012, B1 => n6356, B2 => 
                           n9009, ZN => n1050);
   U2018 : OAI221_X1 port map( B1 => n8955, B2 => n8143, C1 => n6781, C2 => 
                           n8952, A => n1077, ZN => n1074);
   U2019 : AOI22_X1 port map( A1 => n8949, A2 => n8239, B1 => n3321, B2 => 
                           n8946, ZN => n1077);
   U2020 : OAI221_X1 port map( B1 => n8967, B2 => n7983, C1 => n6757, C2 => 
                           n8964, A => n1076, ZN => n1075);
   U2021 : AOI22_X1 port map( A1 => n8961, A2 => n8063, B1 => n8958, B2 => 
                           OUT2_10_port, ZN => n1076);
   U2022 : OAI221_X1 port map( B1 => n8943, B2 => n7801, C1 => n8940, C2 => 
                           n8007, A => n1078, ZN => n1073);
   U2023 : AOI22_X1 port map( A1 => n3404, A2 => n8937, B1 => n3369, B2 => 
                           n8934, ZN => n1078);
   U2024 : OAI221_X1 port map( B1 => n8931, B2 => n7802, C1 => n8928, C2 => 
                           n8039, A => n1079, ZN => n1072);
   U2025 : AOI22_X1 port map( A1 => n3521, A2 => n8925, B1 => n3777, B2 => 
                           n8922, ZN => n1079);
   U2026 : OAI221_X1 port map( B1 => n9018, B2 => n7887, C1 => n9015, C2 => 
                           n8167, A => n1068, ZN => n1067);
   U2027 : AOI22_X1 port map( A1 => n6645, A2 => n9012, B1 => n6357, B2 => 
                           n9009, ZN => n1068);
   U2028 : OAI221_X1 port map( B1 => n8955, B2 => n8144, C1 => n6782, C2 => 
                           n8952, A => n1095, ZN => n1092);
   U2029 : AOI22_X1 port map( A1 => n8949, A2 => n8240, B1 => n3322, B2 => 
                           n8946, ZN => n1095);
   U2030 : OAI221_X1 port map( B1 => n8967, B2 => n7984, C1 => n6758, C2 => 
                           n8964, A => n1094, ZN => n1093);
   U2031 : AOI22_X1 port map( A1 => n8961, A2 => n8064, B1 => n8958, B2 => 
                           OUT2_11_port, ZN => n1094);
   U2032 : OAI221_X1 port map( B1 => n8943, B2 => n7803, C1 => n8940, C2 => 
                           n8008, A => n1096, ZN => n1091);
   U2033 : AOI22_X1 port map( A1 => n3406, A2 => n8937, B1 => n3370, B2 => 
                           n8934, ZN => n1096);
   U2034 : OAI221_X1 port map( B1 => n8931, B2 => n7804, C1 => n8928, C2 => 
                           n8040, A => n1097, ZN => n1090);
   U2035 : AOI22_X1 port map( A1 => n3522, A2 => n8925, B1 => n3778, B2 => 
                           n8922, ZN => n1097);
   U2036 : OAI221_X1 port map( B1 => n9018, B2 => n7888, C1 => n9015, C2 => 
                           n8168, A => n1086, ZN => n1085);
   U2037 : AOI22_X1 port map( A1 => n6646, A2 => n9012, B1 => n6358, B2 => 
                           n9009, ZN => n1086);
   U2038 : OAI221_X1 port map( B1 => n8955, B2 => n8145, C1 => n6783, C2 => 
                           n8952, A => n1113, ZN => n1110);
   U2039 : AOI22_X1 port map( A1 => n8949, A2 => n8241, B1 => n3323, B2 => 
                           n8946, ZN => n1113);
   U2040 : OAI221_X1 port map( B1 => n8967, B2 => n7985, C1 => n6759, C2 => 
                           n8964, A => n1112, ZN => n1111);
   U2041 : AOI22_X1 port map( A1 => n8961, A2 => n8065, B1 => n8958, B2 => 
                           OUT2_12_port, ZN => n1112);
   U2042 : OAI221_X1 port map( B1 => n8943, B2 => n7657, C1 => n8940, C2 => 
                           n8009, A => n1114, ZN => n1109);
   U2043 : AOI22_X1 port map( A1 => n3408, A2 => n8937, B1 => n3371, B2 => 
                           n8934, ZN => n1114);
   U2044 : OAI221_X1 port map( B1 => n8931, B2 => n7658, C1 => n8928, C2 => 
                           n8041, A => n1115, ZN => n1108);
   U2045 : AOI22_X1 port map( A1 => n3523, A2 => n8925, B1 => n3779, B2 => 
                           n8922, ZN => n1115);
   U2046 : OAI221_X1 port map( B1 => n9018, B2 => n7741, C1 => n9015, C2 => 
                           n8169, A => n1104, ZN => n1103);
   U2047 : AOI22_X1 port map( A1 => n6647, A2 => n9012, B1 => n6359, B2 => 
                           n9009, ZN => n1104);
   U2048 : OAI221_X1 port map( B1 => n8955, B2 => n8146, C1 => n6784, C2 => 
                           n8952, A => n1131, ZN => n1128);
   U2049 : AOI22_X1 port map( A1 => n8949, A2 => n8242, B1 => n3324, B2 => 
                           n8946, ZN => n1131);
   U2050 : OAI221_X1 port map( B1 => n8967, B2 => n7986, C1 => n6760, C2 => 
                           n8964, A => n1130, ZN => n1129);
   U2051 : AOI22_X1 port map( A1 => n8961, A2 => n8066, B1 => n8958, B2 => 
                           OUT2_13_port, ZN => n1130);
   U2052 : OAI221_X1 port map( B1 => n8943, B2 => n7659, C1 => n8940, C2 => 
                           n8010, A => n1132, ZN => n1127);
   U2053 : AOI22_X1 port map( A1 => n3410, A2 => n8937, B1 => n3372, B2 => 
                           n8934, ZN => n1132);
   U2054 : OAI221_X1 port map( B1 => n8931, B2 => n7660, C1 => n8928, C2 => 
                           n8042, A => n1133, ZN => n1126);
   U2055 : AOI22_X1 port map( A1 => n3524, A2 => n8925, B1 => n3780, B2 => 
                           n8922, ZN => n1133);
   U2056 : OAI221_X1 port map( B1 => n9018, B2 => n7742, C1 => n9015, C2 => 
                           n8170, A => n1122, ZN => n1121);
   U2057 : AOI22_X1 port map( A1 => n6648, A2 => n9012, B1 => n6360, B2 => 
                           n9009, ZN => n1122);
   U2058 : OAI221_X1 port map( B1 => n8955, B2 => n8147, C1 => n6785, C2 => 
                           n8952, A => n1149, ZN => n1146);
   U2059 : AOI22_X1 port map( A1 => n8949, A2 => n8243, B1 => n3325, B2 => 
                           n8946, ZN => n1149);
   U2060 : OAI221_X1 port map( B1 => n8967, B2 => n7987, C1 => n6761, C2 => 
                           n8964, A => n1148, ZN => n1147);
   U2061 : AOI22_X1 port map( A1 => n8961, A2 => n8067, B1 => n8958, B2 => 
                           OUT2_14_port, ZN => n1148);
   U2062 : OAI221_X1 port map( B1 => n8943, B2 => n7661, C1 => n8940, C2 => 
                           n8011, A => n1150, ZN => n1145);
   U2063 : AOI22_X1 port map( A1 => n3412, A2 => n8937, B1 => n3373, B2 => 
                           n8934, ZN => n1150);
   U2064 : OAI221_X1 port map( B1 => n8931, B2 => n7662, C1 => n8928, C2 => 
                           n8043, A => n1151, ZN => n1144);
   U2065 : AOI22_X1 port map( A1 => n3525, A2 => n8925, B1 => n3781, B2 => 
                           n8922, ZN => n1151);
   U2066 : OAI221_X1 port map( B1 => n9018, B2 => n7743, C1 => n9015, C2 => 
                           n8171, A => n1140, ZN => n1139);
   U2067 : AOI22_X1 port map( A1 => n6649, A2 => n9012, B1 => n6361, B2 => 
                           n9009, ZN => n1140);
   U2068 : OAI221_X1 port map( B1 => n8955, B2 => n8148, C1 => n6786, C2 => 
                           n8952, A => n1167, ZN => n1164);
   U2069 : AOI22_X1 port map( A1 => n8949, A2 => n8244, B1 => n3326, B2 => 
                           n8946, ZN => n1167);
   U2070 : OAI221_X1 port map( B1 => n8967, B2 => n7988, C1 => n6762, C2 => 
                           n8964, A => n1166, ZN => n1165);
   U2071 : AOI22_X1 port map( A1 => n8961, A2 => n8068, B1 => n8958, B2 => 
                           OUT2_15_port, ZN => n1166);
   U2072 : OAI221_X1 port map( B1 => n8943, B2 => n7663, C1 => n8940, C2 => 
                           n8012, A => n1168, ZN => n1163);
   U2073 : AOI22_X1 port map( A1 => n3414, A2 => n8937, B1 => n3374, B2 => 
                           n8934, ZN => n1168);
   U2074 : OAI221_X1 port map( B1 => n8931, B2 => n7664, C1 => n8928, C2 => 
                           n8044, A => n1169, ZN => n1162);
   U2075 : AOI22_X1 port map( A1 => n3526, A2 => n8925, B1 => n3782, B2 => 
                           n8922, ZN => n1169);
   U2076 : OAI221_X1 port map( B1 => n9018, B2 => n7744, C1 => n9015, C2 => 
                           n8172, A => n1158, ZN => n1157);
   U2077 : AOI22_X1 port map( A1 => n6650, A2 => n9012, B1 => n6362, B2 => 
                           n9009, ZN => n1158);
   U2078 : OAI221_X1 port map( B1 => n8955, B2 => n8149, C1 => n6787, C2 => 
                           n8952, A => n1185, ZN => n1182);
   U2079 : AOI22_X1 port map( A1 => n8949, A2 => n8245, B1 => n3327, B2 => 
                           n8946, ZN => n1185);
   U2080 : OAI221_X1 port map( B1 => n8967, B2 => n7989, C1 => n6763, C2 => 
                           n8964, A => n1184, ZN => n1183);
   U2081 : AOI22_X1 port map( A1 => n8961, A2 => n8069, B1 => n8958, B2 => 
                           OUT2_16_port, ZN => n1184);
   U2082 : OAI221_X1 port map( B1 => n8943, B2 => n7665, C1 => n8940, C2 => 
                           n8013, A => n1186, ZN => n1181);
   U2083 : AOI22_X1 port map( A1 => n3416, A2 => n8937, B1 => n3375, B2 => 
                           n8934, ZN => n1186);
   U2084 : OAI221_X1 port map( B1 => n8931, B2 => n7666, C1 => n8928, C2 => 
                           n8045, A => n1187, ZN => n1180);
   U2085 : AOI22_X1 port map( A1 => n3527, A2 => n8925, B1 => n3783, B2 => 
                           n8922, ZN => n1187);
   U2086 : OAI221_X1 port map( B1 => n9018, B2 => n7745, C1 => n9015, C2 => 
                           n8173, A => n1176, ZN => n1175);
   U2087 : AOI22_X1 port map( A1 => n6651, A2 => n9012, B1 => n6363, B2 => 
                           n9009, ZN => n1176);
   U2088 : OAI221_X1 port map( B1 => n8955, B2 => n8150, C1 => n6788, C2 => 
                           n8952, A => n1203, ZN => n1200);
   U2089 : AOI22_X1 port map( A1 => n8949, A2 => n8246, B1 => n3328, B2 => 
                           n8946, ZN => n1203);
   U2090 : OAI221_X1 port map( B1 => n8967, B2 => n7990, C1 => n6764, C2 => 
                           n8964, A => n1202, ZN => n1201);
   U2091 : AOI22_X1 port map( A1 => n8961, A2 => n8070, B1 => n8958, B2 => 
                           OUT2_17_port, ZN => n1202);
   U2092 : OAI221_X1 port map( B1 => n8943, B2 => n7667, C1 => n8940, C2 => 
                           n8014, A => n1204, ZN => n1199);
   U2093 : AOI22_X1 port map( A1 => n3418, A2 => n8937, B1 => n3376, B2 => 
                           n8934, ZN => n1204);
   U2094 : OAI221_X1 port map( B1 => n8931, B2 => n7668, C1 => n8928, C2 => 
                           n8046, A => n1205, ZN => n1198);
   U2095 : AOI22_X1 port map( A1 => n3528, A2 => n8925, B1 => n3784, B2 => 
                           n8922, ZN => n1205);
   U2096 : OAI221_X1 port map( B1 => n9018, B2 => n7746, C1 => n9015, C2 => 
                           n8174, A => n1194, ZN => n1193);
   U2097 : AOI22_X1 port map( A1 => n6652, A2 => n9012, B1 => n6364, B2 => 
                           n9009, ZN => n1194);
   U2098 : OAI221_X1 port map( B1 => n8955, B2 => n8151, C1 => n6789, C2 => 
                           n8952, A => n1221, ZN => n1218);
   U2099 : AOI22_X1 port map( A1 => n8949, A2 => n8247, B1 => n3329, B2 => 
                           n8946, ZN => n1221);
   U2100 : OAI221_X1 port map( B1 => n8967, B2 => n7991, C1 => n6765, C2 => 
                           n8964, A => n1220, ZN => n1219);
   U2101 : AOI22_X1 port map( A1 => n8961, A2 => n8071, B1 => n8958, B2 => 
                           OUT2_18_port, ZN => n1220);
   U2102 : OAI221_X1 port map( B1 => n8943, B2 => n7669, C1 => n8940, C2 => 
                           n8015, A => n1222, ZN => n1217);
   U2103 : AOI22_X1 port map( A1 => n3420, A2 => n8937, B1 => n3377, B2 => 
                           n8934, ZN => n1222);
   U2104 : OAI221_X1 port map( B1 => n8931, B2 => n7670, C1 => n8928, C2 => 
                           n8047, A => n1223, ZN => n1216);
   U2105 : AOI22_X1 port map( A1 => n3529, A2 => n8925, B1 => n3785, B2 => 
                           n8922, ZN => n1223);
   U2106 : OAI221_X1 port map( B1 => n9018, B2 => n7747, C1 => n9015, C2 => 
                           n8175, A => n1212, ZN => n1211);
   U2107 : AOI22_X1 port map( A1 => n6653, A2 => n9012, B1 => n6365, B2 => 
                           n9009, ZN => n1212);
   U2108 : OAI221_X1 port map( B1 => n8955, B2 => n8152, C1 => n6790, C2 => 
                           n8952, A => n1239, ZN => n1236);
   U2109 : AOI22_X1 port map( A1 => n8949, A2 => n8248, B1 => n3330, B2 => 
                           n8946, ZN => n1239);
   U2110 : OAI221_X1 port map( B1 => n8967, B2 => n7992, C1 => n6766, C2 => 
                           n8964, A => n1238, ZN => n1237);
   U2111 : AOI22_X1 port map( A1 => n8961, A2 => n8072, B1 => n8958, B2 => 
                           OUT2_19_port, ZN => n1238);
   U2112 : OAI221_X1 port map( B1 => n8943, B2 => n7671, C1 => n8940, C2 => 
                           n8016, A => n1240, ZN => n1235);
   U2113 : AOI22_X1 port map( A1 => n3422, A2 => n8937, B1 => n3378, B2 => 
                           n8934, ZN => n1240);
   U2114 : OAI221_X1 port map( B1 => n8931, B2 => n7672, C1 => n8928, C2 => 
                           n8048, A => n1241, ZN => n1234);
   U2115 : AOI22_X1 port map( A1 => n3530, A2 => n8925, B1 => n3786, B2 => 
                           n8922, ZN => n1241);
   U2116 : OAI221_X1 port map( B1 => n9018, B2 => n7748, C1 => n9015, C2 => 
                           n8176, A => n1230, ZN => n1229);
   U2117 : AOI22_X1 port map( A1 => n6654, A2 => n9012, B1 => n6366, B2 => 
                           n9009, ZN => n1230);
   U2118 : OAI221_X1 port map( B1 => n8954, B2 => n8153, C1 => n6791, C2 => 
                           n8951, A => n1257, ZN => n1254);
   U2119 : AOI22_X1 port map( A1 => n8948, A2 => n8249, B1 => n3331, B2 => 
                           n8945, ZN => n1257);
   U2120 : OAI221_X1 port map( B1 => n8966, B2 => n7993, C1 => n6767, C2 => 
                           n8963, A => n1256, ZN => n1255);
   U2121 : AOI22_X1 port map( A1 => n8960, A2 => n8073, B1 => n8958, B2 => 
                           OUT2_20_port, ZN => n1256);
   U2122 : OAI221_X1 port map( B1 => n8942, B2 => n7673, C1 => n8939, C2 => 
                           n8017, A => n1258, ZN => n1253);
   U2123 : AOI22_X1 port map( A1 => n3424, A2 => n8936, B1 => n3379, B2 => 
                           n8933, ZN => n1258);
   U2124 : OAI221_X1 port map( B1 => n8930, B2 => n7674, C1 => n8927, C2 => 
                           n8049, A => n1259, ZN => n1252);
   U2125 : AOI22_X1 port map( A1 => n3531, A2 => n8924, B1 => n3787, B2 => 
                           n8921, ZN => n1259);
   U2126 : OAI221_X1 port map( B1 => n9017, B2 => n7749, C1 => n9014, C2 => 
                           n8177, A => n1248, ZN => n1247);
   U2127 : AOI22_X1 port map( A1 => n6655, A2 => n9011, B1 => n6367, B2 => 
                           n9008, ZN => n1248);
   U2128 : OAI221_X1 port map( B1 => n8954, B2 => n8154, C1 => n6792, C2 => 
                           n8951, A => n2299, ZN => n2296);
   U2129 : AOI22_X1 port map( A1 => n8948, A2 => n8250, B1 => n3332, B2 => 
                           n8945, ZN => n2299);
   U2130 : OAI221_X1 port map( B1 => n8966, B2 => n7994, C1 => n6768, C2 => 
                           n8963, A => n2298, ZN => n2297);
   U2131 : AOI22_X1 port map( A1 => n8960, A2 => n8074, B1 => n8959, B2 => 
                           OUT2_21_port, ZN => n2298);
   U2132 : OAI221_X1 port map( B1 => n8942, B2 => n7675, C1 => n8939, C2 => 
                           n8018, A => n2300, ZN => n1271);
   U2133 : AOI22_X1 port map( A1 => n3426, A2 => n8936, B1 => n3380, B2 => 
                           n8933, ZN => n2300);
   U2134 : OAI221_X1 port map( B1 => n8930, B2 => n7676, C1 => n8927, C2 => 
                           n8050, A => n2301, ZN => n1270);
   U2135 : AOI22_X1 port map( A1 => n3532, A2 => n8924, B1 => n3788, B2 => 
                           n8921, ZN => n2301);
   U2136 : OAI221_X1 port map( B1 => n9017, B2 => n7750, C1 => n9014, C2 => 
                           n8178, A => n1266, ZN => n1265);
   U2137 : AOI22_X1 port map( A1 => n6656, A2 => n9011, B1 => n6368, B2 => 
                           n9008, ZN => n1266);
   U2138 : OAI221_X1 port map( B1 => n8954, B2 => n8155, C1 => n6793, C2 => 
                           n8951, A => n2317, ZN => n2314);
   U2139 : AOI22_X1 port map( A1 => n8948, A2 => n8251, B1 => n3333, B2 => 
                           n8945, ZN => n2317);
   U2140 : OAI221_X1 port map( B1 => n8966, B2 => n7995, C1 => n6769, C2 => 
                           n8963, A => n2316, ZN => n2315);
   U2141 : AOI22_X1 port map( A1 => n8960, A2 => n8075, B1 => n8959, B2 => 
                           OUT2_22_port, ZN => n2316);
   U2142 : OAI221_X1 port map( B1 => n8942, B2 => n7677, C1 => n8939, C2 => 
                           n8019, A => n2318, ZN => n2313);
   U2143 : AOI22_X1 port map( A1 => n3428, A2 => n8936, B1 => n3381, B2 => 
                           n8933, ZN => n2318);
   U2144 : OAI221_X1 port map( B1 => n8930, B2 => n7678, C1 => n8927, C2 => 
                           n8051, A => n2319, ZN => n2312);
   U2145 : AOI22_X1 port map( A1 => n3533, A2 => n8924, B1 => n3789, B2 => 
                           n8921, ZN => n2319);
   U2146 : OAI221_X1 port map( B1 => n9017, B2 => n7751, C1 => n9014, C2 => 
                           n8179, A => n2308, ZN => n2307);
   U2147 : AOI22_X1 port map( A1 => n6657, A2 => n9011, B1 => n6369, B2 => 
                           n9008, ZN => n2308);
   U2148 : OAI221_X1 port map( B1 => n8954, B2 => n8156, C1 => n6794, C2 => 
                           n8951, A => n2335, ZN => n2332);
   U2149 : AOI22_X1 port map( A1 => n8948, A2 => n8252, B1 => n3334, B2 => 
                           n8945, ZN => n2335);
   U2150 : OAI221_X1 port map( B1 => n8966, B2 => n7996, C1 => n6770, C2 => 
                           n8963, A => n2334, ZN => n2333);
   U2151 : AOI22_X1 port map( A1 => n8960, A2 => n8076, B1 => n8959, B2 => 
                           OUT2_23_port, ZN => n2334);
   U2152 : OAI221_X1 port map( B1 => n8942, B2 => n7679, C1 => n8939, C2 => 
                           n8020, A => n2336, ZN => n2331);
   U2153 : AOI22_X1 port map( A1 => n3430, A2 => n8936, B1 => n3382, B2 => 
                           n8933, ZN => n2336);
   U2154 : OAI221_X1 port map( B1 => n8930, B2 => n7680, C1 => n8927, C2 => 
                           n8052, A => n2337, ZN => n2330);
   U2155 : AOI22_X1 port map( A1 => n3534, A2 => n8924, B1 => n3790, B2 => 
                           n8921, ZN => n2337);
   U2156 : OAI221_X1 port map( B1 => n9017, B2 => n7752, C1 => n9014, C2 => 
                           n8180, A => n2326, ZN => n2325);
   U2157 : AOI22_X1 port map( A1 => n6658, A2 => n9011, B1 => n6370, B2 => 
                           n9008, ZN => n2326);
   U2158 : OAI221_X1 port map( B1 => n8954, B2 => n7869, C1 => n6739, C2 => 
                           n8951, A => n2353, ZN => n2350);
   U2159 : AOI22_X1 port map( A1 => n8948, A2 => n8253, B1 => n3263, B2 => 
                           n8945, ZN => n2353);
   U2160 : OAI221_X1 port map( B1 => n8966, B2 => n7805, C1 => n6731, C2 => 
                           n8963, A => n2352, ZN => n2351);
   U2161 : AOI22_X1 port map( A1 => n8960, A2 => n8077, B1 => n8959, B2 => 
                           OUT2_24_port, ZN => n2352);
   U2162 : OAI221_X1 port map( B1 => n8942, B2 => n7806, C1 => n8939, C2 => 
                           n8021, A => n2354, ZN => n2349);
   U2163 : AOI22_X1 port map( A1 => n3432, A2 => n8936, B1 => n3279, B2 => 
                           n8933, ZN => n2354);
   U2164 : OAI221_X1 port map( B1 => n8930, B2 => n7681, C1 => n8927, C2 => 
                           n7821, A => n2355, ZN => n2348);
   U2165 : AOI22_X1 port map( A1 => n3535, A2 => n8924, B1 => n3567, B2 => 
                           n8921, ZN => n2355);
   U2166 : OAI221_X1 port map( B1 => n9017, B2 => n7753, C1 => n9014, C2 => 
                           n7901, A => n2344, ZN => n2343);
   U2167 : AOI22_X1 port map( A1 => n6659, A2 => n9011, B1 => n6371, B2 => 
                           n9008, ZN => n2344);
   U2168 : OAI221_X1 port map( B1 => n8954, B2 => n7870, C1 => n6740, C2 => 
                           n8951, A => n2371, ZN => n2368);
   U2169 : AOI22_X1 port map( A1 => n8948, A2 => n8254, B1 => n3264, B2 => 
                           n8945, ZN => n2371);
   U2170 : OAI221_X1 port map( B1 => n8966, B2 => n7807, C1 => n6732, C2 => 
                           n8963, A => n2370, ZN => n2369);
   U2171 : AOI22_X1 port map( A1 => n8960, A2 => n8078, B1 => n8959, B2 => 
                           OUT2_25_port, ZN => n2370);
   U2172 : OAI221_X1 port map( B1 => n8942, B2 => n7808, C1 => n8939, C2 => 
                           n8022, A => n2372, ZN => n2367);
   U2173 : AOI22_X1 port map( A1 => n3434, A2 => n8936, B1 => n3280, B2 => 
                           n8933, ZN => n2372);
   U2174 : OAI221_X1 port map( B1 => n8930, B2 => n7682, C1 => n8927, C2 => 
                           n7822, A => n2373, ZN => n2366);
   U2175 : AOI22_X1 port map( A1 => n3536, A2 => n8924, B1 => n3568, B2 => 
                           n8921, ZN => n2373);
   U2176 : OAI221_X1 port map( B1 => n9017, B2 => n7754, C1 => n9014, C2 => 
                           n7902, A => n2362, ZN => n2361);
   U2177 : AOI22_X1 port map( A1 => n6660, A2 => n9011, B1 => n6372, B2 => 
                           n9008, ZN => n2362);
   U2178 : OAI221_X1 port map( B1 => n8954, B2 => n7871, C1 => n6741, C2 => 
                           n8951, A => n2389, ZN => n2386);
   U2179 : AOI22_X1 port map( A1 => n8948, A2 => n8255, B1 => n3265, B2 => 
                           n8945, ZN => n2389);
   U2180 : OAI221_X1 port map( B1 => n8966, B2 => n7809, C1 => n6733, C2 => 
                           n8963, A => n2388, ZN => n2387);
   U2181 : AOI22_X1 port map( A1 => n8960, A2 => n8079, B1 => n8959, B2 => 
                           OUT2_26_port, ZN => n2388);
   U2182 : OAI221_X1 port map( B1 => n8942, B2 => n7810, C1 => n8939, C2 => 
                           n8023, A => n2390, ZN => n2385);
   U2183 : AOI22_X1 port map( A1 => n3436, A2 => n8936, B1 => n3281, B2 => 
                           n8933, ZN => n2390);
   U2184 : OAI221_X1 port map( B1 => n8930, B2 => n7683, C1 => n8927, C2 => 
                           n7823, A => n2391, ZN => n2384);
   U2185 : AOI22_X1 port map( A1 => n3537, A2 => n8924, B1 => n3569, B2 => 
                           n8921, ZN => n2391);
   U2186 : OAI221_X1 port map( B1 => n9017, B2 => n7755, C1 => n9014, C2 => 
                           n7903, A => n2380, ZN => n2379);
   U2187 : AOI22_X1 port map( A1 => n6661, A2 => n9011, B1 => n6373, B2 => 
                           n9008, ZN => n2380);
   U2188 : OAI221_X1 port map( B1 => n8954, B2 => n7872, C1 => n6742, C2 => 
                           n8951, A => n2407, ZN => n2404);
   U2189 : AOI22_X1 port map( A1 => n8948, A2 => n8256, B1 => n3266, B2 => 
                           n8945, ZN => n2407);
   U2190 : OAI221_X1 port map( B1 => n8966, B2 => n7811, C1 => n6734, C2 => 
                           n8963, A => n2406, ZN => n2405);
   U2191 : AOI22_X1 port map( A1 => n8960, A2 => n8080, B1 => n8959, B2 => 
                           OUT2_27_port, ZN => n2406);
   U2192 : OAI221_X1 port map( B1 => n8942, B2 => n7812, C1 => n8939, C2 => 
                           n8024, A => n2408, ZN => n2403);
   U2193 : AOI22_X1 port map( A1 => n3438, A2 => n8936, B1 => n3282, B2 => 
                           n8933, ZN => n2408);
   U2194 : OAI221_X1 port map( B1 => n8930, B2 => n7684, C1 => n8927, C2 => 
                           n7824, A => n2409, ZN => n2402);
   U2195 : AOI22_X1 port map( A1 => n3538, A2 => n8924, B1 => n3570, B2 => 
                           n8921, ZN => n2409);
   U2196 : OAI221_X1 port map( B1 => n9017, B2 => n7756, C1 => n9014, C2 => 
                           n7904, A => n2398, ZN => n2397);
   U2197 : AOI22_X1 port map( A1 => n6662, A2 => n9011, B1 => n6374, B2 => 
                           n9008, ZN => n2398);
   U2198 : OAI221_X1 port map( B1 => n8954, B2 => n7873, C1 => n6743, C2 => 
                           n8951, A => n2425, ZN => n2422);
   U2199 : AOI22_X1 port map( A1 => n8948, A2 => n8257, B1 => n3267, B2 => 
                           n8945, ZN => n2425);
   U2200 : OAI221_X1 port map( B1 => n8966, B2 => n7813, C1 => n6735, C2 => 
                           n8963, A => n2424, ZN => n2423);
   U2201 : AOI22_X1 port map( A1 => n8960, A2 => n8081, B1 => n8959, B2 => 
                           OUT2_28_port, ZN => n2424);
   U2202 : OAI221_X1 port map( B1 => n8942, B2 => n7814, C1 => n8939, C2 => 
                           n8025, A => n2426, ZN => n2421);
   U2203 : AOI22_X1 port map( A1 => n3440, A2 => n8936, B1 => n3283, B2 => 
                           n8933, ZN => n2426);
   U2204 : OAI221_X1 port map( B1 => n8930, B2 => n7685, C1 => n8927, C2 => 
                           n7825, A => n2427, ZN => n2420);
   U2205 : AOI22_X1 port map( A1 => n3539, A2 => n8924, B1 => n3571, B2 => 
                           n8921, ZN => n2427);
   U2206 : OAI221_X1 port map( B1 => n9017, B2 => n7757, C1 => n9014, C2 => 
                           n7905, A => n2416, ZN => n2415);
   U2207 : AOI22_X1 port map( A1 => n6663, A2 => n9011, B1 => n6375, B2 => 
                           n9008, ZN => n2416);
   U2208 : OAI221_X1 port map( B1 => n8954, B2 => n7874, C1 => n6744, C2 => 
                           n8951, A => n2443, ZN => n2440);
   U2209 : AOI22_X1 port map( A1 => n8948, A2 => n8258, B1 => n3268, B2 => 
                           n8945, ZN => n2443);
   U2210 : OAI221_X1 port map( B1 => n8966, B2 => n7815, C1 => n6736, C2 => 
                           n8963, A => n2442, ZN => n2441);
   U2211 : AOI22_X1 port map( A1 => n8960, A2 => n8082, B1 => n8959, B2 => 
                           OUT2_29_port, ZN => n2442);
   U2212 : OAI221_X1 port map( B1 => n8942, B2 => n7816, C1 => n8939, C2 => 
                           n8026, A => n2444, ZN => n2439);
   U2213 : AOI22_X1 port map( A1 => n3442, A2 => n8936, B1 => n3284, B2 => 
                           n8933, ZN => n2444);
   U2214 : OAI221_X1 port map( B1 => n8930, B2 => n7686, C1 => n8927, C2 => 
                           n7826, A => n2445, ZN => n2438);
   U2215 : AOI22_X1 port map( A1 => n3540, A2 => n8924, B1 => n3572, B2 => 
                           n8921, ZN => n2445);
   U2216 : OAI221_X1 port map( B1 => n9017, B2 => n7758, C1 => n9014, C2 => 
                           n7906, A => n2434, ZN => n2433);
   U2217 : AOI22_X1 port map( A1 => n6664, A2 => n9011, B1 => n6376, B2 => 
                           n9008, ZN => n2434);
   U2218 : OAI221_X1 port map( B1 => n8954, B2 => n7875, C1 => n6745, C2 => 
                           n8951, A => n2461, ZN => n2458);
   U2219 : AOI22_X1 port map( A1 => n8948, A2 => n8259, B1 => n3269, B2 => 
                           n8945, ZN => n2461);
   U2220 : OAI221_X1 port map( B1 => n8966, B2 => n7817, C1 => n6737, C2 => 
                           n8963, A => n2460, ZN => n2459);
   U2221 : AOI22_X1 port map( A1 => n8960, A2 => n8083, B1 => n8959, B2 => 
                           OUT2_30_port, ZN => n2460);
   U2222 : OAI221_X1 port map( B1 => n8942, B2 => n7818, C1 => n8939, C2 => 
                           n8027, A => n2462, ZN => n2457);
   U2223 : AOI22_X1 port map( A1 => n3444, A2 => n8936, B1 => n3285, B2 => 
                           n8933, ZN => n2462);
   U2224 : OAI221_X1 port map( B1 => n8930, B2 => n7687, C1 => n8927, C2 => 
                           n7827, A => n2463, ZN => n2456);
   U2225 : AOI22_X1 port map( A1 => n3541, A2 => n8924, B1 => n3573, B2 => 
                           n8921, ZN => n2463);
   U2226 : OAI221_X1 port map( B1 => n9017, B2 => n7759, C1 => n9014, C2 => 
                           n7907, A => n2452, ZN => n2451);
   U2227 : AOI22_X1 port map( A1 => n6665, A2 => n9011, B1 => n6377, B2 => 
                           n9008, ZN => n2452);
   U2228 : OAI221_X1 port map( B1 => n8954, B2 => n7876, C1 => n6746, C2 => 
                           n8951, A => n2490, ZN => n2486);
   U2229 : AOI22_X1 port map( A1 => n8948, A2 => n8260, B1 => n3270, B2 => 
                           n8945, ZN => n2490);
   U2230 : OAI221_X1 port map( B1 => n8966, B2 => n7819, C1 => n6738, C2 => 
                           n8963, A => n2488, ZN => n2487);
   U2231 : AOI22_X1 port map( A1 => n8960, A2 => n8084, B1 => n8957, B2 => 
                           OUT2_31_port, ZN => n2488);
   U2232 : OAI221_X1 port map( B1 => n8942, B2 => n7820, C1 => n8939, C2 => 
                           n8028, A => n2492, ZN => n2485);
   U2233 : AOI22_X1 port map( A1 => n3446, A2 => n8936, B1 => n3286, B2 => 
                           n8933, ZN => n2492);
   U2234 : OAI221_X1 port map( B1 => n8930, B2 => n7688, C1 => n8927, C2 => 
                           n7828, A => n2493, ZN => n2484);
   U2235 : AOI22_X1 port map( A1 => n3542, A2 => n8924, B1 => n3574, B2 => 
                           n8921, ZN => n2493);
   U2236 : OAI221_X1 port map( B1 => n9017, B2 => n7760, C1 => n9014, C2 => 
                           n7908, A => n2470, ZN => n2469);
   U2237 : AOI22_X1 port map( A1 => n6666, A2 => n9011, B1 => n6378, B2 => 
                           n9008, ZN => n2470);
   U2238 : OAI221_X1 port map( B1 => n6835, B2 => n8908, C1 => n8205, C2 => 
                           n8905, A => n2509, ZN => n2500);
   U2239 : AOI22_X1 port map( A1 => n8902, A2 => n3335, B1 => n8897, B2 => 
                           n8261, ZN => n2509);
   U2240 : OAI221_X1 port map( B1 => n6836, B2 => n8908, C1 => n8206, C2 => 
                           n8905, A => n2554, ZN => n2551);
   U2241 : AOI22_X1 port map( A1 => n8902, A2 => n3336, B1 => n8897, B2 => 
                           n8262, ZN => n2554);
   U2242 : OAI221_X1 port map( B1 => n6837, B2 => n8908, C1 => n8207, C2 => 
                           n8905, A => n2572, ZN => n2569);
   U2243 : AOI22_X1 port map( A1 => n8902, A2 => n3337, B1 => n8897, B2 => 
                           n8263, ZN => n2572);
   U2244 : OAI221_X1 port map( B1 => n6838, B2 => n8908, C1 => n8208, C2 => 
                           n8905, A => n2590, ZN => n2587);
   U2245 : AOI22_X1 port map( A1 => n8902, A2 => n3338, B1 => n8897, B2 => 
                           n8264, ZN => n2590);
   U2246 : OAI221_X1 port map( B1 => n6839, B2 => n8908, C1 => n8209, C2 => 
                           n8905, A => n2608, ZN => n2605);
   U2247 : AOI22_X1 port map( A1 => n8902, A2 => n3339, B1 => n8897, B2 => 
                           n8265, ZN => n2608);
   U2248 : OAI221_X1 port map( B1 => n6840, B2 => n8908, C1 => n8210, C2 => 
                           n8905, A => n2626, ZN => n2623);
   U2249 : AOI22_X1 port map( A1 => n8902, A2 => n3340, B1 => n8897, B2 => 
                           n8266, ZN => n2626);
   U2250 : OAI221_X1 port map( B1 => n6841, B2 => n8908, C1 => n8211, C2 => 
                           n8905, A => n2644, ZN => n2641);
   U2251 : AOI22_X1 port map( A1 => n8902, A2 => n3341, B1 => n8897, B2 => 
                           n8267, ZN => n2644);
   U2252 : OAI221_X1 port map( B1 => n6842, B2 => n8908, C1 => n8212, C2 => 
                           n8905, A => n2662, ZN => n2659);
   U2253 : AOI22_X1 port map( A1 => n8902, A2 => n3342, B1 => n8897, B2 => 
                           n8268, ZN => n2662);
   U2254 : OAI221_X1 port map( B1 => n6843, B2 => n8907, C1 => n8213, C2 => 
                           n8904, A => n2680, ZN => n2677);
   U2255 : AOI22_X1 port map( A1 => n8901, A2 => n3343, B1 => n8897, B2 => 
                           n8269, ZN => n2680);
   U2256 : OAI221_X1 port map( B1 => n6844, B2 => n8907, C1 => n8214, C2 => 
                           n8904, A => n2698, ZN => n2695);
   U2257 : AOI22_X1 port map( A1 => n8901, A2 => n3344, B1 => n8897, B2 => 
                           n8270, ZN => n2698);
   U2258 : OAI221_X1 port map( B1 => n6845, B2 => n8907, C1 => n8215, C2 => 
                           n8904, A => n2716, ZN => n2713);
   U2259 : AOI22_X1 port map( A1 => n8901, A2 => n3345, B1 => n8897, B2 => 
                           n8271, ZN => n2716);
   U2260 : OAI221_X1 port map( B1 => n6846, B2 => n8907, C1 => n8216, C2 => 
                           n8904, A => n2734, ZN => n2731);
   U2261 : AOI22_X1 port map( A1 => n8901, A2 => n3346, B1 => n8897, B2 => 
                           n8272, ZN => n2734);
   U2262 : OAI221_X1 port map( B1 => n6847, B2 => n8907, C1 => n8217, C2 => 
                           n8904, A => n2752, ZN => n2749);
   U2263 : AOI22_X1 port map( A1 => n8901, A2 => n3347, B1 => n8898, B2 => 
                           n8273, ZN => n2752);
   U2264 : OAI221_X1 port map( B1 => n6848, B2 => n8907, C1 => n8218, C2 => 
                           n8904, A => n2770, ZN => n2767);
   U2265 : AOI22_X1 port map( A1 => n8901, A2 => n3348, B1 => n8898, B2 => 
                           n8274, ZN => n2770);
   U2266 : OAI221_X1 port map( B1 => n6849, B2 => n8907, C1 => n8219, C2 => 
                           n8904, A => n2788, ZN => n2785);
   U2267 : AOI22_X1 port map( A1 => n8901, A2 => n3349, B1 => n8898, B2 => 
                           n8275, ZN => n2788);
   U2268 : OAI221_X1 port map( B1 => n6850, B2 => n8907, C1 => n8220, C2 => 
                           n8904, A => n2806, ZN => n2803);
   U2269 : AOI22_X1 port map( A1 => n8901, A2 => n3350, B1 => n8898, B2 => 
                           n8276, ZN => n2806);
   U2270 : OAI221_X1 port map( B1 => n6851, B2 => n8907, C1 => n8221, C2 => 
                           n8904, A => n2824, ZN => n2821);
   U2271 : AOI22_X1 port map( A1 => n8901, A2 => n3351, B1 => n8898, B2 => 
                           n8277, ZN => n2824);
   U2272 : OAI221_X1 port map( B1 => n6852, B2 => n8907, C1 => n8222, C2 => 
                           n8904, A => n2842, ZN => n2839);
   U2273 : AOI22_X1 port map( A1 => n8901, A2 => n3352, B1 => n8898, B2 => 
                           n8278, ZN => n2842);
   U2274 : OAI221_X1 port map( B1 => n6853, B2 => n8907, C1 => n8223, C2 => 
                           n8904, A => n2860, ZN => n2857);
   U2275 : AOI22_X1 port map( A1 => n8901, A2 => n3353, B1 => n8898, B2 => 
                           n8279, ZN => n2860);
   U2276 : OAI221_X1 port map( B1 => n6854, B2 => n8907, C1 => n8224, C2 => 
                           n8904, A => n2878, ZN => n2875);
   U2277 : AOI22_X1 port map( A1 => n8901, A2 => n3354, B1 => n8898, B2 => 
                           n8280, ZN => n2878);
   U2278 : OAI221_X1 port map( B1 => n6855, B2 => n8906, C1 => n8225, C2 => 
                           n8903, A => n2896, ZN => n2893);
   U2279 : AOI22_X1 port map( A1 => n8900, A2 => n3355, B1 => n8898, B2 => 
                           n8281, ZN => n2896);
   U2280 : OAI221_X1 port map( B1 => n6856, B2 => n8906, C1 => n8226, C2 => 
                           n8903, A => n2914, ZN => n2911);
   U2281 : AOI22_X1 port map( A1 => n8900, A2 => n3356, B1 => n8898, B2 => 
                           n8282, ZN => n2914);
   U2282 : OAI221_X1 port map( B1 => n6857, B2 => n8906, C1 => n8227, C2 => 
                           n8903, A => n2932, ZN => n2929);
   U2283 : AOI22_X1 port map( A1 => n8900, A2 => n3357, B1 => n8898, B2 => 
                           n8283, ZN => n2932);
   U2284 : OAI221_X1 port map( B1 => n6858, B2 => n8906, C1 => n8228, C2 => 
                           n8903, A => n2950, ZN => n2947);
   U2285 : AOI22_X1 port map( A1 => n8900, A2 => n3358, B1 => n8898, B2 => 
                           n8284, ZN => n2950);
   U2286 : OAI221_X1 port map( B1 => n6803, B2 => n8906, C1 => n7917, C2 => 
                           n8903, A => n2968, ZN => n2965);
   U2287 : AOI22_X1 port map( A1 => n8900, A2 => n3271, B1 => n8899, B2 => 
                           n8285, ZN => n2968);
   U2288 : OAI221_X1 port map( B1 => n6804, B2 => n8906, C1 => n7918, C2 => 
                           n8903, A => n2986, ZN => n2983);
   U2289 : AOI22_X1 port map( A1 => n8900, A2 => n3272, B1 => n8899, B2 => 
                           n8286, ZN => n2986);
   U2290 : OAI221_X1 port map( B1 => n6805, B2 => n8906, C1 => n7919, C2 => 
                           n8903, A => n3004, ZN => n3001);
   U2291 : AOI22_X1 port map( A1 => n8900, A2 => n3273, B1 => n8899, B2 => 
                           n8287, ZN => n3004);
   U2292 : OAI221_X1 port map( B1 => n6806, B2 => n8906, C1 => n7920, C2 => 
                           n8903, A => n3022, ZN => n3019);
   U2293 : AOI22_X1 port map( A1 => n8900, A2 => n3274, B1 => n8899, B2 => 
                           n8288, ZN => n3022);
   U2294 : OAI221_X1 port map( B1 => n6807, B2 => n8906, C1 => n7921, C2 => 
                           n8903, A => n3040, ZN => n3037);
   U2295 : AOI22_X1 port map( A1 => n8900, A2 => n3275, B1 => n8899, B2 => 
                           n8289, ZN => n3040);
   U2296 : OAI221_X1 port map( B1 => n6808, B2 => n8906, C1 => n7922, C2 => 
                           n8903, A => n3058, ZN => n3055);
   U2297 : AOI22_X1 port map( A1 => n8900, A2 => n3276, B1 => n8899, B2 => 
                           n8290, ZN => n3058);
   U2298 : OAI221_X1 port map( B1 => n6809, B2 => n8906, C1 => n7923, C2 => 
                           n8903, A => n3076, ZN => n3073);
   U2299 : AOI22_X1 port map( A1 => n8900, A2 => n3277, B1 => n8899, B2 => 
                           n8291, ZN => n3076);
   U2300 : OAI221_X1 port map( B1 => n6810, B2 => n8906, C1 => n7924, C2 => 
                           n8903, A => n3098, ZN => n3091);
   U2301 : AOI22_X1 port map( A1 => n8900, A2 => n3278, B1 => n8899, B2 => 
                           n8292, ZN => n3098);
   U2302 : OAI22_X1 port map( A1 => n8673, A2 => n8717, B1 => n6835, B2 => 
                           n8672, ZN => n2104);
   U2303 : OAI22_X1 port map( A1 => n8673, A2 => n8720, B1 => n6836, B2 => 
                           n8672, ZN => n2105);
   U2304 : OAI22_X1 port map( A1 => n8673, A2 => n8723, B1 => n6837, B2 => 
                           n8672, ZN => n2106);
   U2305 : OAI22_X1 port map( A1 => n8673, A2 => n8726, B1 => n6838, B2 => 
                           n8672, ZN => n2107);
   U2306 : OAI22_X1 port map( A1 => n8673, A2 => n8729, B1 => n6839, B2 => 
                           n8672, ZN => n2108);
   U2307 : OAI22_X1 port map( A1 => n8674, A2 => n8732, B1 => n6840, B2 => 
                           n8672, ZN => n2109);
   U2308 : OAI22_X1 port map( A1 => n8674, A2 => n8735, B1 => n6841, B2 => 
                           n8672, ZN => n2110);
   U2309 : OAI22_X1 port map( A1 => n8674, A2 => n8738, B1 => n6842, B2 => 
                           n8672, ZN => n2111);
   U2310 : OAI22_X1 port map( A1 => n8674, A2 => n8741, B1 => n6843, B2 => 
                           n8672, ZN => n2112);
   U2311 : OAI22_X1 port map( A1 => n8674, A2 => n8744, B1 => n6844, B2 => 
                           n8672, ZN => n2113);
   U2312 : OAI22_X1 port map( A1 => n8675, A2 => n8747, B1 => n6845, B2 => 
                           n8672, ZN => n2114);
   U2313 : OAI22_X1 port map( A1 => n8675, A2 => n8750, B1 => n6846, B2 => 
                           n8672, ZN => n2115);
   U2314 : OAI22_X1 port map( A1 => n8675, A2 => n8753, B1 => n6847, B2 => 
                           n3158, ZN => n2116);
   U2315 : OAI22_X1 port map( A1 => n8675, A2 => n8756, B1 => n6848, B2 => 
                           n3158, ZN => n2117);
   U2316 : OAI22_X1 port map( A1 => n8675, A2 => n8759, B1 => n6849, B2 => 
                           n3158, ZN => n2118);
   U2317 : OAI22_X1 port map( A1 => n8676, A2 => n8762, B1 => n6850, B2 => 
                           n8672, ZN => n2119);
   U2318 : OAI22_X1 port map( A1 => n8676, A2 => n8765, B1 => n6851, B2 => 
                           n8672, ZN => n2120);
   U2319 : OAI22_X1 port map( A1 => n8676, A2 => n8768, B1 => n6852, B2 => 
                           n8672, ZN => n2121);
   U2320 : OAI22_X1 port map( A1 => n8676, A2 => n8771, B1 => n6853, B2 => 
                           n8672, ZN => n2122);
   U2321 : OAI22_X1 port map( A1 => n8676, A2 => n8774, B1 => n6854, B2 => 
                           n8672, ZN => n2123);
   U2322 : OAI22_X1 port map( A1 => n8677, A2 => n8777, B1 => n6855, B2 => 
                           n8672, ZN => n2124);
   U2323 : OAI22_X1 port map( A1 => n8677, A2 => n8780, B1 => n6856, B2 => 
                           n8672, ZN => n2125);
   U2324 : OAI22_X1 port map( A1 => n8677, A2 => n8783, B1 => n6857, B2 => 
                           n8672, ZN => n2126);
   U2325 : OAI22_X1 port map( A1 => n8677, A2 => n8786, B1 => n6858, B2 => 
                           n8672, ZN => n2127);
   U2326 : OAI22_X1 port map( A1 => n8448, A2 => n8719, B1 => n6627, B2 => 
                           n8447, ZN => n1304);
   U2327 : OAI22_X1 port map( A1 => n8448, A2 => n8722, B1 => n6628, B2 => 
                           n8447, ZN => n1305);
   U2328 : OAI22_X1 port map( A1 => n8448, A2 => n8725, B1 => n6629, B2 => 
                           n8447, ZN => n1306);
   U2329 : OAI22_X1 port map( A1 => n8448, A2 => n8728, B1 => n6630, B2 => 
                           n8447, ZN => n1307);
   U2330 : OAI22_X1 port map( A1 => n8448, A2 => n8731, B1 => n6631, B2 => 
                           n8447, ZN => n1308);
   U2331 : OAI22_X1 port map( A1 => n8449, A2 => n8734, B1 => n6632, B2 => 
                           n8447, ZN => n1309);
   U2332 : OAI22_X1 port map( A1 => n8449, A2 => n8737, B1 => n6633, B2 => 
                           n8447, ZN => n1310);
   U2333 : OAI22_X1 port map( A1 => n8449, A2 => n8740, B1 => n6634, B2 => 
                           n8447, ZN => n1311);
   U2334 : OAI22_X1 port map( A1 => n8449, A2 => n8743, B1 => n6603, B2 => 
                           n8447, ZN => n1312);
   U2335 : OAI22_X1 port map( A1 => n8449, A2 => n8746, B1 => n6604, B2 => 
                           n8447, ZN => n1313);
   U2336 : OAI22_X1 port map( A1 => n8450, A2 => n8749, B1 => n6605, B2 => 
                           n8447, ZN => n1314);
   U2337 : OAI22_X1 port map( A1 => n8450, A2 => n8752, B1 => n6606, B2 => 
                           n8447, ZN => n1315);
   U2338 : OAI22_X1 port map( A1 => n8450, A2 => n8755, B1 => n6607, B2 => 
                           n3189, ZN => n1316);
   U2339 : OAI22_X1 port map( A1 => n8450, A2 => n8758, B1 => n6608, B2 => 
                           n3189, ZN => n1317);
   U2340 : OAI22_X1 port map( A1 => n8450, A2 => n8761, B1 => n6609, B2 => 
                           n3189, ZN => n1318);
   U2341 : OAI22_X1 port map( A1 => n8451, A2 => n8764, B1 => n6610, B2 => 
                           n8447, ZN => n1319);
   U2342 : OAI22_X1 port map( A1 => n8451, A2 => n8767, B1 => n6611, B2 => 
                           n8447, ZN => n1320);
   U2343 : OAI22_X1 port map( A1 => n8451, A2 => n8770, B1 => n6612, B2 => 
                           n8447, ZN => n1321);
   U2344 : OAI22_X1 port map( A1 => n8451, A2 => n8773, B1 => n6613, B2 => 
                           n8447, ZN => n1322);
   U2345 : OAI22_X1 port map( A1 => n8451, A2 => n8776, B1 => n6614, B2 => 
                           n8447, ZN => n1323);
   U2346 : OAI22_X1 port map( A1 => n8452, A2 => n8779, B1 => n6615, B2 => 
                           n8447, ZN => n1324);
   U2347 : OAI22_X1 port map( A1 => n8452, A2 => n8782, B1 => n6616, B2 => 
                           n8447, ZN => n1325);
   U2348 : OAI22_X1 port map( A1 => n8452, A2 => n8785, B1 => n6617, B2 => 
                           n8447, ZN => n1326);
   U2349 : OAI22_X1 port map( A1 => n8452, A2 => n8788, B1 => n6618, B2 => 
                           n8447, ZN => n1327);
   U2350 : OAI22_X1 port map( A1 => n8457, A2 => n8719, B1 => n8341, B2 => 
                           n8456, ZN => n1336);
   U2351 : OAI22_X1 port map( A1 => n8457, A2 => n8722, B1 => n8342, B2 => 
                           n8456, ZN => n1337);
   U2352 : OAI22_X1 port map( A1 => n8457, A2 => n8725, B1 => n8343, B2 => 
                           n8456, ZN => n1338);
   U2353 : OAI22_X1 port map( A1 => n8457, A2 => n8728, B1 => n8344, B2 => 
                           n8456, ZN => n1339);
   U2354 : OAI22_X1 port map( A1 => n8457, A2 => n8731, B1 => n8345, B2 => 
                           n8456, ZN => n1340);
   U2355 : OAI22_X1 port map( A1 => n8458, A2 => n8734, B1 => n8346, B2 => 
                           n8456, ZN => n1341);
   U2356 : OAI22_X1 port map( A1 => n8458, A2 => n8737, B1 => n8347, B2 => 
                           n8456, ZN => n1342);
   U2357 : OAI22_X1 port map( A1 => n8458, A2 => n8740, B1 => n8348, B2 => 
                           n8456, ZN => n1343);
   U2358 : OAI22_X1 port map( A1 => n8458, A2 => n8743, B1 => n8349, B2 => 
                           n8456, ZN => n1344);
   U2359 : OAI22_X1 port map( A1 => n8458, A2 => n8746, B1 => n8350, B2 => 
                           n8456, ZN => n1345);
   U2360 : OAI22_X1 port map( A1 => n8459, A2 => n8749, B1 => n8351, B2 => 
                           n8456, ZN => n1346);
   U2361 : OAI22_X1 port map( A1 => n8459, A2 => n8752, B1 => n8352, B2 => 
                           n8456, ZN => n1347);
   U2362 : OAI22_X1 port map( A1 => n8459, A2 => n8755, B1 => n8353, B2 => 
                           n3188, ZN => n1348);
   U2363 : OAI22_X1 port map( A1 => n8459, A2 => n8758, B1 => n8354, B2 => 
                           n3188, ZN => n1349);
   U2364 : OAI22_X1 port map( A1 => n8459, A2 => n8761, B1 => n8355, B2 => 
                           n3188, ZN => n1350);
   U2365 : OAI22_X1 port map( A1 => n8460, A2 => n8764, B1 => n8356, B2 => 
                           n8456, ZN => n1351);
   U2366 : OAI22_X1 port map( A1 => n8460, A2 => n8767, B1 => n8357, B2 => 
                           n8456, ZN => n1352);
   U2367 : OAI22_X1 port map( A1 => n8460, A2 => n8770, B1 => n8358, B2 => 
                           n8456, ZN => n1353);
   U2368 : OAI22_X1 port map( A1 => n8460, A2 => n8773, B1 => n8359, B2 => 
                           n8456, ZN => n1354);
   U2369 : OAI22_X1 port map( A1 => n8460, A2 => n8776, B1 => n8360, B2 => 
                           n8456, ZN => n1355);
   U2370 : OAI22_X1 port map( A1 => n8461, A2 => n8779, B1 => n8361, B2 => 
                           n8456, ZN => n1356);
   U2371 : OAI22_X1 port map( A1 => n8461, A2 => n8782, B1 => n8362, B2 => 
                           n8456, ZN => n1357);
   U2372 : OAI22_X1 port map( A1 => n8461, A2 => n8785, B1 => n8363, B2 => 
                           n8456, ZN => n1358);
   U2373 : OAI22_X1 port map( A1 => n8461, A2 => n8788, B1 => n8364, B2 => 
                           n8456, ZN => n1359);
   U2374 : OAI22_X1 port map( A1 => n8466, A2 => n8719, B1 => n8365, B2 => 
                           n8465, ZN => n1368);
   U2375 : OAI22_X1 port map( A1 => n8466, A2 => n8722, B1 => n8366, B2 => 
                           n8465, ZN => n1369);
   U2376 : OAI22_X1 port map( A1 => n8466, A2 => n8725, B1 => n8367, B2 => 
                           n8465, ZN => n1370);
   U2377 : OAI22_X1 port map( A1 => n8466, A2 => n8728, B1 => n8368, B2 => 
                           n8465, ZN => n1371);
   U2378 : OAI22_X1 port map( A1 => n8466, A2 => n8731, B1 => n8369, B2 => 
                           n8465, ZN => n1372);
   U2379 : OAI22_X1 port map( A1 => n8467, A2 => n8734, B1 => n8370, B2 => 
                           n8465, ZN => n1373);
   U2380 : OAI22_X1 port map( A1 => n8467, A2 => n8737, B1 => n8371, B2 => 
                           n8465, ZN => n1374);
   U2381 : OAI22_X1 port map( A1 => n8467, A2 => n8740, B1 => n8372, B2 => 
                           n8465, ZN => n1375);
   U2382 : OAI22_X1 port map( A1 => n8467, A2 => n8743, B1 => n8373, B2 => 
                           n8465, ZN => n1376);
   U2383 : OAI22_X1 port map( A1 => n8467, A2 => n8746, B1 => n8374, B2 => 
                           n8465, ZN => n1377);
   U2384 : OAI22_X1 port map( A1 => n8468, A2 => n8749, B1 => n8375, B2 => 
                           n8465, ZN => n1378);
   U2385 : OAI22_X1 port map( A1 => n8468, A2 => n8752, B1 => n8376, B2 => 
                           n8465, ZN => n1379);
   U2386 : OAI22_X1 port map( A1 => n8468, A2 => n8755, B1 => n8377, B2 => 
                           n3187, ZN => n1380);
   U2387 : OAI22_X1 port map( A1 => n8468, A2 => n8758, B1 => n8378, B2 => 
                           n3187, ZN => n1381);
   U2388 : OAI22_X1 port map( A1 => n8468, A2 => n8761, B1 => n8379, B2 => 
                           n3187, ZN => n1382);
   U2389 : OAI22_X1 port map( A1 => n8469, A2 => n8764, B1 => n8380, B2 => 
                           n8465, ZN => n1383);
   U2390 : OAI22_X1 port map( A1 => n8469, A2 => n8767, B1 => n8381, B2 => 
                           n8465, ZN => n1384);
   U2391 : OAI22_X1 port map( A1 => n8469, A2 => n8770, B1 => n8382, B2 => 
                           n8465, ZN => n1385);
   U2392 : OAI22_X1 port map( A1 => n8469, A2 => n8773, B1 => n8383, B2 => 
                           n8465, ZN => n1386);
   U2393 : OAI22_X1 port map( A1 => n8469, A2 => n8776, B1 => n8384, B2 => 
                           n8465, ZN => n1387);
   U2394 : OAI22_X1 port map( A1 => n8470, A2 => n8779, B1 => n8385, B2 => 
                           n8465, ZN => n1388);
   U2395 : OAI22_X1 port map( A1 => n8470, A2 => n8782, B1 => n8386, B2 => 
                           n8465, ZN => n1389);
   U2396 : OAI22_X1 port map( A1 => n8470, A2 => n8785, B1 => n8387, B2 => 
                           n8465, ZN => n1390);
   U2397 : OAI22_X1 port map( A1 => n8470, A2 => n8788, B1 => n8388, B2 => 
                           n8465, ZN => n1391);
   U2398 : OAI22_X1 port map( A1 => n8484, A2 => n8719, B1 => n6683, B2 => 
                           n8483, ZN => n1432);
   U2399 : OAI22_X1 port map( A1 => n8484, A2 => n8722, B1 => n6684, B2 => 
                           n8483, ZN => n1433);
   U2400 : OAI22_X1 port map( A1 => n8484, A2 => n8725, B1 => n6685, B2 => 
                           n8483, ZN => n1434);
   U2401 : OAI22_X1 port map( A1 => n8484, A2 => n8728, B1 => n6686, B2 => 
                           n8483, ZN => n1435);
   U2402 : OAI22_X1 port map( A1 => n8484, A2 => n8731, B1 => n6687, B2 => 
                           n8483, ZN => n1436);
   U2403 : OAI22_X1 port map( A1 => n8485, A2 => n8734, B1 => n6688, B2 => 
                           n8483, ZN => n1437);
   U2404 : OAI22_X1 port map( A1 => n8485, A2 => n8737, B1 => n6689, B2 => 
                           n8483, ZN => n1438);
   U2405 : OAI22_X1 port map( A1 => n8485, A2 => n8740, B1 => n6690, B2 => 
                           n8483, ZN => n1439);
   U2406 : OAI22_X1 port map( A1 => n8485, A2 => n8743, B1 => n6691, B2 => 
                           n8483, ZN => n1440);
   U2407 : OAI22_X1 port map( A1 => n8485, A2 => n8746, B1 => n6692, B2 => 
                           n8483, ZN => n1441);
   U2408 : OAI22_X1 port map( A1 => n8486, A2 => n8749, B1 => n6693, B2 => 
                           n8483, ZN => n1442);
   U2409 : OAI22_X1 port map( A1 => n8486, A2 => n8752, B1 => n6694, B2 => 
                           n8483, ZN => n1443);
   U2410 : OAI22_X1 port map( A1 => n8486, A2 => n8755, B1 => n6695, B2 => 
                           n3185, ZN => n1444);
   U2411 : OAI22_X1 port map( A1 => n8486, A2 => n8758, B1 => n6696, B2 => 
                           n3185, ZN => n1445);
   U2412 : OAI22_X1 port map( A1 => n8486, A2 => n8761, B1 => n6697, B2 => 
                           n3185, ZN => n1446);
   U2413 : OAI22_X1 port map( A1 => n8487, A2 => n8764, B1 => n6698, B2 => 
                           n8483, ZN => n1447);
   U2414 : OAI22_X1 port map( A1 => n8487, A2 => n8767, B1 => n6699, B2 => 
                           n8483, ZN => n1448);
   U2415 : OAI22_X1 port map( A1 => n8487, A2 => n8770, B1 => n6700, B2 => 
                           n8483, ZN => n1449);
   U2416 : OAI22_X1 port map( A1 => n8487, A2 => n8773, B1 => n6701, B2 => 
                           n8483, ZN => n1450);
   U2417 : OAI22_X1 port map( A1 => n8487, A2 => n8776, B1 => n6702, B2 => 
                           n8483, ZN => n1451);
   U2418 : OAI22_X1 port map( A1 => n8488, A2 => n8779, B1 => n6703, B2 => 
                           n8483, ZN => n1452);
   U2419 : OAI22_X1 port map( A1 => n8488, A2 => n8782, B1 => n6704, B2 => 
                           n8483, ZN => n1453);
   U2420 : OAI22_X1 port map( A1 => n8488, A2 => n8785, B1 => n6705, B2 => 
                           n8483, ZN => n1454);
   U2421 : OAI22_X1 port map( A1 => n8488, A2 => n8788, B1 => n6706, B2 => 
                           n8483, ZN => n1455);
   U2422 : OAI22_X1 port map( A1 => n8502, A2 => n8719, B1 => n6875, B2 => 
                           n8501, ZN => n1496);
   U2423 : OAI22_X1 port map( A1 => n8502, A2 => n8722, B1 => n6876, B2 => 
                           n8501, ZN => n1497);
   U2424 : OAI22_X1 port map( A1 => n8502, A2 => n8725, B1 => n6877, B2 => 
                           n8501, ZN => n1498);
   U2425 : OAI22_X1 port map( A1 => n8502, A2 => n8728, B1 => n6878, B2 => 
                           n8501, ZN => n1499);
   U2426 : OAI22_X1 port map( A1 => n8502, A2 => n8731, B1 => n6879, B2 => 
                           n8501, ZN => n1500);
   U2427 : OAI22_X1 port map( A1 => n8503, A2 => n8734, B1 => n6880, B2 => 
                           n8501, ZN => n1501);
   U2428 : OAI22_X1 port map( A1 => n8503, A2 => n8737, B1 => n6881, B2 => 
                           n8501, ZN => n1502);
   U2429 : OAI22_X1 port map( A1 => n8503, A2 => n8740, B1 => n6882, B2 => 
                           n8501, ZN => n1503);
   U2430 : OAI22_X1 port map( A1 => n8503, A2 => n8743, B1 => n6883, B2 => 
                           n8501, ZN => n1504);
   U2431 : OAI22_X1 port map( A1 => n8503, A2 => n8746, B1 => n6884, B2 => 
                           n8501, ZN => n1505);
   U2432 : OAI22_X1 port map( A1 => n8504, A2 => n8749, B1 => n6885, B2 => 
                           n8501, ZN => n1506);
   U2433 : OAI22_X1 port map( A1 => n8504, A2 => n8752, B1 => n6886, B2 => 
                           n8501, ZN => n1507);
   U2434 : OAI22_X1 port map( A1 => n8504, A2 => n8755, B1 => n6887, B2 => 
                           n3182, ZN => n1508);
   U2435 : OAI22_X1 port map( A1 => n8504, A2 => n8758, B1 => n6888, B2 => 
                           n3182, ZN => n1509);
   U2436 : OAI22_X1 port map( A1 => n8504, A2 => n8761, B1 => n6889, B2 => 
                           n3182, ZN => n1510);
   U2437 : OAI22_X1 port map( A1 => n8505, A2 => n8764, B1 => n6890, B2 => 
                           n8501, ZN => n1511);
   U2438 : OAI22_X1 port map( A1 => n8505, A2 => n8767, B1 => n6891, B2 => 
                           n8501, ZN => n1512);
   U2439 : OAI22_X1 port map( A1 => n8505, A2 => n8770, B1 => n6892, B2 => 
                           n8501, ZN => n1513);
   U2440 : OAI22_X1 port map( A1 => n8505, A2 => n8773, B1 => n6893, B2 => 
                           n8501, ZN => n1514);
   U2441 : OAI22_X1 port map( A1 => n8505, A2 => n8776, B1 => n6894, B2 => 
                           n8501, ZN => n1515);
   U2442 : OAI22_X1 port map( A1 => n8506, A2 => n8779, B1 => n6895, B2 => 
                           n8501, ZN => n1516);
   U2443 : OAI22_X1 port map( A1 => n8506, A2 => n8782, B1 => n6896, B2 => 
                           n8501, ZN => n1517);
   U2444 : OAI22_X1 port map( A1 => n8506, A2 => n8785, B1 => n6897, B2 => 
                           n8501, ZN => n1518);
   U2445 : OAI22_X1 port map( A1 => n8506, A2 => n8788, B1 => n6898, B2 => 
                           n8501, ZN => n1519);
   U2446 : OAI22_X1 port map( A1 => n8511, A2 => n8718, B1 => n8293, B2 => 
                           n8510, ZN => n1528);
   U2447 : OAI22_X1 port map( A1 => n8511, A2 => n8721, B1 => n8294, B2 => 
                           n8510, ZN => n1529);
   U2448 : OAI22_X1 port map( A1 => n8511, A2 => n8724, B1 => n8295, B2 => 
                           n8510, ZN => n1530);
   U2449 : OAI22_X1 port map( A1 => n8511, A2 => n8727, B1 => n8296, B2 => 
                           n8510, ZN => n1531);
   U2450 : OAI22_X1 port map( A1 => n8511, A2 => n8730, B1 => n8297, B2 => 
                           n8510, ZN => n1532);
   U2451 : OAI22_X1 port map( A1 => n8512, A2 => n8733, B1 => n8298, B2 => 
                           n8510, ZN => n1533);
   U2452 : OAI22_X1 port map( A1 => n8512, A2 => n8736, B1 => n8299, B2 => 
                           n8510, ZN => n1534);
   U2453 : OAI22_X1 port map( A1 => n8512, A2 => n8739, B1 => n8300, B2 => 
                           n8510, ZN => n1535);
   U2454 : OAI22_X1 port map( A1 => n8512, A2 => n8742, B1 => n8301, B2 => 
                           n8510, ZN => n1536);
   U2455 : OAI22_X1 port map( A1 => n8512, A2 => n8745, B1 => n8302, B2 => 
                           n8510, ZN => n1537);
   U2456 : OAI22_X1 port map( A1 => n8513, A2 => n8748, B1 => n8303, B2 => 
                           n8510, ZN => n1538);
   U2457 : OAI22_X1 port map( A1 => n8513, A2 => n8751, B1 => n8304, B2 => 
                           n8510, ZN => n1539);
   U2458 : OAI22_X1 port map( A1 => n8513, A2 => n8754, B1 => n8305, B2 => 
                           n3181, ZN => n1540);
   U2459 : OAI22_X1 port map( A1 => n8513, A2 => n8757, B1 => n8306, B2 => 
                           n3181, ZN => n1541);
   U2460 : OAI22_X1 port map( A1 => n8513, A2 => n8760, B1 => n8307, B2 => 
                           n3181, ZN => n1542);
   U2461 : OAI22_X1 port map( A1 => n8514, A2 => n8763, B1 => n8308, B2 => 
                           n8510, ZN => n1543);
   U2462 : OAI22_X1 port map( A1 => n8514, A2 => n8766, B1 => n8309, B2 => 
                           n8510, ZN => n1544);
   U2463 : OAI22_X1 port map( A1 => n8514, A2 => n8769, B1 => n8310, B2 => 
                           n8510, ZN => n1545);
   U2464 : OAI22_X1 port map( A1 => n8514, A2 => n8772, B1 => n8311, B2 => 
                           n8510, ZN => n1546);
   U2465 : OAI22_X1 port map( A1 => n8514, A2 => n8775, B1 => n8312, B2 => 
                           n8510, ZN => n1547);
   U2466 : OAI22_X1 port map( A1 => n8515, A2 => n8778, B1 => n8313, B2 => 
                           n8510, ZN => n1548);
   U2467 : OAI22_X1 port map( A1 => n8515, A2 => n8781, B1 => n8314, B2 => 
                           n8510, ZN => n1549);
   U2468 : OAI22_X1 port map( A1 => n8515, A2 => n8784, B1 => n8315, B2 => 
                           n8510, ZN => n1550);
   U2469 : OAI22_X1 port map( A1 => n8515, A2 => n8787, B1 => n8316, B2 => 
                           n8510, ZN => n1551);
   U2470 : OAI22_X1 port map( A1 => n8529, A2 => n8718, B1 => n6339, B2 => 
                           n8528, ZN => n1592);
   U2471 : OAI22_X1 port map( A1 => n8529, A2 => n8721, B1 => n6340, B2 => 
                           n8528, ZN => n1593);
   U2472 : OAI22_X1 port map( A1 => n8529, A2 => n8724, B1 => n6341, B2 => 
                           n8528, ZN => n1594);
   U2473 : OAI22_X1 port map( A1 => n8529, A2 => n8727, B1 => n6342, B2 => 
                           n8528, ZN => n1595);
   U2474 : OAI22_X1 port map( A1 => n8529, A2 => n8730, B1 => n6343, B2 => 
                           n8528, ZN => n1596);
   U2475 : OAI22_X1 port map( A1 => n8530, A2 => n8733, B1 => n6344, B2 => 
                           n8528, ZN => n1597);
   U2476 : OAI22_X1 port map( A1 => n8530, A2 => n8736, B1 => n6345, B2 => 
                           n8528, ZN => n1598);
   U2477 : OAI22_X1 port map( A1 => n8530, A2 => n8739, B1 => n6346, B2 => 
                           n8528, ZN => n1599);
   U2478 : OAI22_X1 port map( A1 => n8530, A2 => n8742, B1 => n6315, B2 => 
                           n8528, ZN => n1600);
   U2479 : OAI22_X1 port map( A1 => n8530, A2 => n8745, B1 => n6316, B2 => 
                           n8528, ZN => n1601);
   U2480 : OAI22_X1 port map( A1 => n8531, A2 => n8748, B1 => n6317, B2 => 
                           n8528, ZN => n1602);
   U2481 : OAI22_X1 port map( A1 => n8531, A2 => n8751, B1 => n6318, B2 => 
                           n8528, ZN => n1603);
   U2482 : OAI22_X1 port map( A1 => n8531, A2 => n8754, B1 => n6319, B2 => 
                           n3179, ZN => n1604);
   U2483 : OAI22_X1 port map( A1 => n8531, A2 => n8757, B1 => n6320, B2 => 
                           n3179, ZN => n1605);
   U2484 : OAI22_X1 port map( A1 => n8531, A2 => n8760, B1 => n6321, B2 => 
                           n3179, ZN => n1606);
   U2485 : OAI22_X1 port map( A1 => n8532, A2 => n8763, B1 => n6322, B2 => 
                           n8528, ZN => n1607);
   U2486 : OAI22_X1 port map( A1 => n8532, A2 => n8766, B1 => n6323, B2 => 
                           n8528, ZN => n1608);
   U2487 : OAI22_X1 port map( A1 => n8532, A2 => n8769, B1 => n6324, B2 => 
                           n8528, ZN => n1609);
   U2488 : OAI22_X1 port map( A1 => n8532, A2 => n8772, B1 => n6325, B2 => 
                           n8528, ZN => n1610);
   U2489 : OAI22_X1 port map( A1 => n8532, A2 => n8775, B1 => n6326, B2 => 
                           n8528, ZN => n1611);
   U2490 : OAI22_X1 port map( A1 => n8533, A2 => n8778, B1 => n6327, B2 => 
                           n8528, ZN => n1612);
   U2491 : OAI22_X1 port map( A1 => n8533, A2 => n8781, B1 => n6328, B2 => 
                           n8528, ZN => n1613);
   U2492 : OAI22_X1 port map( A1 => n8533, A2 => n8784, B1 => n6329, B2 => 
                           n8528, ZN => n1614);
   U2493 : OAI22_X1 port map( A1 => n8533, A2 => n8787, B1 => n6330, B2 => 
                           n8528, ZN => n1615);
   U2494 : OAI22_X1 port map( A1 => n8547, A2 => n8718, B1 => n8317, B2 => 
                           n8546, ZN => n1656);
   U2495 : OAI22_X1 port map( A1 => n8547, A2 => n8721, B1 => n8318, B2 => 
                           n8546, ZN => n1657);
   U2496 : OAI22_X1 port map( A1 => n8547, A2 => n8724, B1 => n8319, B2 => 
                           n8546, ZN => n1658);
   U2497 : OAI22_X1 port map( A1 => n8547, A2 => n8727, B1 => n8320, B2 => 
                           n8546, ZN => n1659);
   U2498 : OAI22_X1 port map( A1 => n8547, A2 => n8730, B1 => n8321, B2 => 
                           n8546, ZN => n1660);
   U2499 : OAI22_X1 port map( A1 => n8548, A2 => n8733, B1 => n8322, B2 => 
                           n8546, ZN => n1661);
   U2500 : OAI22_X1 port map( A1 => n8548, A2 => n8736, B1 => n8323, B2 => 
                           n8546, ZN => n1662);
   U2501 : OAI22_X1 port map( A1 => n8548, A2 => n8739, B1 => n8324, B2 => 
                           n8546, ZN => n1663);
   U2502 : OAI22_X1 port map( A1 => n8548, A2 => n8742, B1 => n8325, B2 => 
                           n8546, ZN => n1664);
   U2503 : OAI22_X1 port map( A1 => n8548, A2 => n8745, B1 => n8326, B2 => 
                           n8546, ZN => n1665);
   U2504 : OAI22_X1 port map( A1 => n8549, A2 => n8748, B1 => n8327, B2 => 
                           n8546, ZN => n1666);
   U2505 : OAI22_X1 port map( A1 => n8549, A2 => n8751, B1 => n8328, B2 => 
                           n8546, ZN => n1667);
   U2506 : OAI22_X1 port map( A1 => n8549, A2 => n8754, B1 => n8329, B2 => 
                           n3177, ZN => n1668);
   U2507 : OAI22_X1 port map( A1 => n8549, A2 => n8757, B1 => n8330, B2 => 
                           n3177, ZN => n1669);
   U2508 : OAI22_X1 port map( A1 => n8549, A2 => n8760, B1 => n8331, B2 => 
                           n3177, ZN => n1670);
   U2509 : OAI22_X1 port map( A1 => n8550, A2 => n8763, B1 => n8332, B2 => 
                           n8546, ZN => n1671);
   U2510 : OAI22_X1 port map( A1 => n8550, A2 => n8766, B1 => n8333, B2 => 
                           n8546, ZN => n1672);
   U2511 : OAI22_X1 port map( A1 => n8550, A2 => n8769, B1 => n8334, B2 => 
                           n8546, ZN => n1673);
   U2512 : OAI22_X1 port map( A1 => n8550, A2 => n8772, B1 => n8335, B2 => 
                           n8546, ZN => n1674);
   U2513 : OAI22_X1 port map( A1 => n8550, A2 => n8775, B1 => n8336, B2 => 
                           n8546, ZN => n1675);
   U2514 : OAI22_X1 port map( A1 => n8551, A2 => n8778, B1 => n8337, B2 => 
                           n8546, ZN => n1676);
   U2515 : OAI22_X1 port map( A1 => n8551, A2 => n8781, B1 => n8338, B2 => 
                           n8546, ZN => n1677);
   U2516 : OAI22_X1 port map( A1 => n8551, A2 => n8784, B1 => n8339, B2 => 
                           n8546, ZN => n1678);
   U2517 : OAI22_X1 port map( A1 => n8551, A2 => n8787, B1 => n8340, B2 => 
                           n8546, ZN => n1679);
   U2518 : OAI22_X1 port map( A1 => n8556, A2 => n8718, B1 => n6707, B2 => 
                           n8555, ZN => n1688);
   U2519 : OAI22_X1 port map( A1 => n8556, A2 => n8721, B1 => n6708, B2 => 
                           n8555, ZN => n1689);
   U2520 : OAI22_X1 port map( A1 => n8556, A2 => n8724, B1 => n6709, B2 => 
                           n8555, ZN => n1690);
   U2521 : OAI22_X1 port map( A1 => n8556, A2 => n8727, B1 => n6710, B2 => 
                           n8555, ZN => n1691);
   U2522 : OAI22_X1 port map( A1 => n8556, A2 => n8730, B1 => n6711, B2 => 
                           n8555, ZN => n1692);
   U2523 : OAI22_X1 port map( A1 => n8557, A2 => n8733, B1 => n6712, B2 => 
                           n8555, ZN => n1693);
   U2524 : OAI22_X1 port map( A1 => n8557, A2 => n8736, B1 => n6713, B2 => 
                           n8555, ZN => n1694);
   U2525 : OAI22_X1 port map( A1 => n8557, A2 => n8739, B1 => n6714, B2 => 
                           n8555, ZN => n1695);
   U2526 : OAI22_X1 port map( A1 => n8557, A2 => n8742, B1 => n6715, B2 => 
                           n8555, ZN => n1696);
   U2527 : OAI22_X1 port map( A1 => n8557, A2 => n8745, B1 => n6716, B2 => 
                           n8555, ZN => n1697);
   U2528 : OAI22_X1 port map( A1 => n8558, A2 => n8748, B1 => n6717, B2 => 
                           n8555, ZN => n1698);
   U2529 : OAI22_X1 port map( A1 => n8558, A2 => n8751, B1 => n6718, B2 => 
                           n8555, ZN => n1699);
   U2530 : OAI22_X1 port map( A1 => n8558, A2 => n8754, B1 => n6719, B2 => 
                           n3176, ZN => n1700);
   U2531 : OAI22_X1 port map( A1 => n8558, A2 => n8757, B1 => n6720, B2 => 
                           n3176, ZN => n1701);
   U2532 : OAI22_X1 port map( A1 => n8558, A2 => n8760, B1 => n6721, B2 => 
                           n3176, ZN => n1702);
   U2533 : OAI22_X1 port map( A1 => n8559, A2 => n8763, B1 => n6722, B2 => 
                           n8555, ZN => n1703);
   U2534 : OAI22_X1 port map( A1 => n8559, A2 => n8766, B1 => n6723, B2 => 
                           n8555, ZN => n1704);
   U2535 : OAI22_X1 port map( A1 => n8559, A2 => n8769, B1 => n6724, B2 => 
                           n8555, ZN => n1705);
   U2536 : OAI22_X1 port map( A1 => n8559, A2 => n8772, B1 => n6725, B2 => 
                           n8555, ZN => n1706);
   U2537 : OAI22_X1 port map( A1 => n8559, A2 => n8775, B1 => n6726, B2 => 
                           n8555, ZN => n1707);
   U2538 : OAI22_X1 port map( A1 => n8560, A2 => n8778, B1 => n6727, B2 => 
                           n8555, ZN => n1708);
   U2539 : OAI22_X1 port map( A1 => n8560, A2 => n8781, B1 => n6728, B2 => 
                           n8555, ZN => n1709);
   U2540 : OAI22_X1 port map( A1 => n8560, A2 => n8784, B1 => n6729, B2 => 
                           n8555, ZN => n1710);
   U2541 : OAI22_X1 port map( A1 => n8560, A2 => n8787, B1 => n6730, B2 => 
                           n8555, ZN => n1711);
   U2542 : OAI22_X1 port map( A1 => n8592, A2 => n8718, B1 => n6811, B2 => 
                           n8591, ZN => n1816);
   U2543 : OAI22_X1 port map( A1 => n8592, A2 => n8721, B1 => n6812, B2 => 
                           n8591, ZN => n1817);
   U2544 : OAI22_X1 port map( A1 => n8592, A2 => n8724, B1 => n6813, B2 => 
                           n8591, ZN => n1818);
   U2545 : OAI22_X1 port map( A1 => n8592, A2 => n8727, B1 => n6814, B2 => 
                           n8591, ZN => n1819);
   U2546 : OAI22_X1 port map( A1 => n8592, A2 => n8730, B1 => n6815, B2 => 
                           n8591, ZN => n1820);
   U2547 : OAI22_X1 port map( A1 => n8593, A2 => n8733, B1 => n6816, B2 => 
                           n8591, ZN => n1821);
   U2548 : OAI22_X1 port map( A1 => n8593, A2 => n8736, B1 => n6817, B2 => 
                           n8591, ZN => n1822);
   U2549 : OAI22_X1 port map( A1 => n8593, A2 => n8739, B1 => n6818, B2 => 
                           n8591, ZN => n1823);
   U2550 : OAI22_X1 port map( A1 => n8593, A2 => n8742, B1 => n6819, B2 => 
                           n8591, ZN => n1824);
   U2551 : OAI22_X1 port map( A1 => n8593, A2 => n8745, B1 => n6820, B2 => 
                           n8591, ZN => n1825);
   U2552 : OAI22_X1 port map( A1 => n8594, A2 => n8748, B1 => n6821, B2 => 
                           n8591, ZN => n1826);
   U2553 : OAI22_X1 port map( A1 => n8594, A2 => n8751, B1 => n6822, B2 => 
                           n8591, ZN => n1827);
   U2554 : OAI22_X1 port map( A1 => n8594, A2 => n8754, B1 => n6823, B2 => 
                           n3171, ZN => n1828);
   U2555 : OAI22_X1 port map( A1 => n8594, A2 => n8757, B1 => n6824, B2 => 
                           n3171, ZN => n1829);
   U2556 : OAI22_X1 port map( A1 => n8594, A2 => n8760, B1 => n6825, B2 => 
                           n3171, ZN => n1830);
   U2557 : OAI22_X1 port map( A1 => n8595, A2 => n8763, B1 => n6826, B2 => 
                           n8591, ZN => n1831);
   U2558 : OAI22_X1 port map( A1 => n8595, A2 => n8766, B1 => n6827, B2 => 
                           n8591, ZN => n1832);
   U2559 : OAI22_X1 port map( A1 => n8595, A2 => n8769, B1 => n6828, B2 => 
                           n8591, ZN => n1833);
   U2560 : OAI22_X1 port map( A1 => n8595, A2 => n8772, B1 => n6829, B2 => 
                           n8591, ZN => n1834);
   U2561 : OAI22_X1 port map( A1 => n8595, A2 => n8775, B1 => n6830, B2 => 
                           n8591, ZN => n1835);
   U2562 : OAI22_X1 port map( A1 => n8596, A2 => n8778, B1 => n6831, B2 => 
                           n8591, ZN => n1836);
   U2563 : OAI22_X1 port map( A1 => n8596, A2 => n8781, B1 => n6832, B2 => 
                           n8591, ZN => n1837);
   U2564 : OAI22_X1 port map( A1 => n8596, A2 => n8784, B1 => n6833, B2 => 
                           n8591, ZN => n1838);
   U2565 : OAI22_X1 port map( A1 => n8596, A2 => n8787, B1 => n6834, B2 => 
                           n8591, ZN => n1839);
   U2566 : OAI22_X1 port map( A1 => n8601, A2 => n8718, B1 => n6747, B2 => 
                           n8600, ZN => n1848);
   U2567 : OAI22_X1 port map( A1 => n8601, A2 => n8721, B1 => n6748, B2 => 
                           n8600, ZN => n1849);
   U2568 : OAI22_X1 port map( A1 => n8601, A2 => n8724, B1 => n6749, B2 => 
                           n8600, ZN => n1850);
   U2569 : OAI22_X1 port map( A1 => n8601, A2 => n8727, B1 => n6750, B2 => 
                           n8600, ZN => n1851);
   U2570 : OAI22_X1 port map( A1 => n8601, A2 => n8730, B1 => n6751, B2 => 
                           n8600, ZN => n1852);
   U2571 : OAI22_X1 port map( A1 => n8602, A2 => n8733, B1 => n6752, B2 => 
                           n8600, ZN => n1853);
   U2572 : OAI22_X1 port map( A1 => n8602, A2 => n8736, B1 => n6753, B2 => 
                           n8600, ZN => n1854);
   U2573 : OAI22_X1 port map( A1 => n8602, A2 => n8739, B1 => n6754, B2 => 
                           n8600, ZN => n1855);
   U2574 : OAI22_X1 port map( A1 => n8602, A2 => n8742, B1 => n6755, B2 => 
                           n8600, ZN => n1856);
   U2575 : OAI22_X1 port map( A1 => n8602, A2 => n8745, B1 => n6756, B2 => 
                           n8600, ZN => n1857);
   U2576 : OAI22_X1 port map( A1 => n8603, A2 => n8748, B1 => n6757, B2 => 
                           n8600, ZN => n1858);
   U2577 : OAI22_X1 port map( A1 => n8603, A2 => n8751, B1 => n6758, B2 => 
                           n8600, ZN => n1859);
   U2578 : OAI22_X1 port map( A1 => n8603, A2 => n8754, B1 => n6759, B2 => 
                           n3170, ZN => n1860);
   U2579 : OAI22_X1 port map( A1 => n8603, A2 => n8757, B1 => n6760, B2 => 
                           n3170, ZN => n1861);
   U2580 : OAI22_X1 port map( A1 => n8603, A2 => n8760, B1 => n6761, B2 => 
                           n3170, ZN => n1862);
   U2581 : OAI22_X1 port map( A1 => n8604, A2 => n8763, B1 => n6762, B2 => 
                           n8600, ZN => n1863);
   U2582 : OAI22_X1 port map( A1 => n8604, A2 => n8766, B1 => n6763, B2 => 
                           n8600, ZN => n1864);
   U2583 : OAI22_X1 port map( A1 => n8604, A2 => n8769, B1 => n6764, B2 => 
                           n8600, ZN => n1865);
   U2584 : OAI22_X1 port map( A1 => n8604, A2 => n8772, B1 => n6765, B2 => 
                           n8600, ZN => n1866);
   U2585 : OAI22_X1 port map( A1 => n8604, A2 => n8775, B1 => n6766, B2 => 
                           n8600, ZN => n1867);
   U2586 : OAI22_X1 port map( A1 => n8605, A2 => n8778, B1 => n6767, B2 => 
                           n8600, ZN => n1868);
   U2587 : OAI22_X1 port map( A1 => n8605, A2 => n8781, B1 => n6768, B2 => 
                           n8600, ZN => n1869);
   U2588 : OAI22_X1 port map( A1 => n8605, A2 => n8784, B1 => n6769, B2 => 
                           n8600, ZN => n1870);
   U2589 : OAI22_X1 port map( A1 => n8605, A2 => n8787, B1 => n6770, B2 => 
                           n8600, ZN => n1871);
   U2590 : OAI22_X1 port map( A1 => n8610, A2 => n8718, B1 => n6771, B2 => 
                           n8609, ZN => n1880);
   U2591 : OAI22_X1 port map( A1 => n8610, A2 => n8721, B1 => n6772, B2 => 
                           n8609, ZN => n1881);
   U2592 : OAI22_X1 port map( A1 => n8610, A2 => n8724, B1 => n6773, B2 => 
                           n8609, ZN => n1882);
   U2593 : OAI22_X1 port map( A1 => n8610, A2 => n8727, B1 => n6774, B2 => 
                           n8609, ZN => n1883);
   U2594 : OAI22_X1 port map( A1 => n8610, A2 => n8730, B1 => n6775, B2 => 
                           n8609, ZN => n1884);
   U2595 : OAI22_X1 port map( A1 => n8611, A2 => n8733, B1 => n6776, B2 => 
                           n8609, ZN => n1885);
   U2596 : OAI22_X1 port map( A1 => n8611, A2 => n8736, B1 => n6777, B2 => 
                           n8609, ZN => n1886);
   U2597 : OAI22_X1 port map( A1 => n8611, A2 => n8739, B1 => n6778, B2 => 
                           n8609, ZN => n1887);
   U2598 : OAI22_X1 port map( A1 => n8611, A2 => n8742, B1 => n6779, B2 => 
                           n8609, ZN => n1888);
   U2599 : OAI22_X1 port map( A1 => n8611, A2 => n8745, B1 => n6780, B2 => 
                           n8609, ZN => n1889);
   U2600 : OAI22_X1 port map( A1 => n8612, A2 => n8748, B1 => n6781, B2 => 
                           n8609, ZN => n1890);
   U2601 : OAI22_X1 port map( A1 => n8612, A2 => n8751, B1 => n6782, B2 => 
                           n8609, ZN => n1891);
   U2602 : OAI22_X1 port map( A1 => n8612, A2 => n8754, B1 => n6783, B2 => 
                           n3169, ZN => n1892);
   U2603 : OAI22_X1 port map( A1 => n8612, A2 => n8757, B1 => n6784, B2 => 
                           n3169, ZN => n1893);
   U2604 : OAI22_X1 port map( A1 => n8612, A2 => n8760, B1 => n6785, B2 => 
                           n3169, ZN => n1894);
   U2605 : OAI22_X1 port map( A1 => n8613, A2 => n8763, B1 => n6786, B2 => 
                           n8609, ZN => n1895);
   U2606 : OAI22_X1 port map( A1 => n8613, A2 => n8766, B1 => n6787, B2 => 
                           n8609, ZN => n1896);
   U2607 : OAI22_X1 port map( A1 => n8613, A2 => n8769, B1 => n6788, B2 => 
                           n8609, ZN => n1897);
   U2608 : OAI22_X1 port map( A1 => n8613, A2 => n8772, B1 => n6789, B2 => 
                           n8609, ZN => n1898);
   U2609 : OAI22_X1 port map( A1 => n8613, A2 => n8775, B1 => n6790, B2 => 
                           n8609, ZN => n1899);
   U2610 : OAI22_X1 port map( A1 => n8614, A2 => n8778, B1 => n6791, B2 => 
                           n8609, ZN => n1900);
   U2611 : OAI22_X1 port map( A1 => n8614, A2 => n8781, B1 => n6792, B2 => 
                           n8609, ZN => n1901);
   U2612 : OAI22_X1 port map( A1 => n8614, A2 => n8784, B1 => n6793, B2 => 
                           n8609, ZN => n1902);
   U2613 : OAI22_X1 port map( A1 => n8614, A2 => n8787, B1 => n6794, B2 => 
                           n8609, ZN => n1903);
   U2614 : OAI22_X1 port map( A1 => n8619, A2 => n8717, B1 => n8389, B2 => 
                           n8618, ZN => n1912);
   U2615 : OAI22_X1 port map( A1 => n8619, A2 => n8720, B1 => n8390, B2 => 
                           n8618, ZN => n1913);
   U2616 : OAI22_X1 port map( A1 => n8619, A2 => n8723, B1 => n8391, B2 => 
                           n8618, ZN => n1914);
   U2617 : OAI22_X1 port map( A1 => n8619, A2 => n8726, B1 => n8392, B2 => 
                           n8618, ZN => n1915);
   U2618 : OAI22_X1 port map( A1 => n8619, A2 => n8729, B1 => n8393, B2 => 
                           n8618, ZN => n1916);
   U2619 : OAI22_X1 port map( A1 => n8620, A2 => n8732, B1 => n8394, B2 => 
                           n8618, ZN => n1917);
   U2620 : OAI22_X1 port map( A1 => n8620, A2 => n8735, B1 => n8395, B2 => 
                           n8618, ZN => n1918);
   U2621 : OAI22_X1 port map( A1 => n8620, A2 => n8738, B1 => n8396, B2 => 
                           n8618, ZN => n1919);
   U2622 : OAI22_X1 port map( A1 => n8620, A2 => n8741, B1 => n8397, B2 => 
                           n8618, ZN => n1920);
   U2623 : OAI22_X1 port map( A1 => n8620, A2 => n8744, B1 => n8398, B2 => 
                           n8618, ZN => n1921);
   U2624 : OAI22_X1 port map( A1 => n8621, A2 => n8747, B1 => n8399, B2 => 
                           n8618, ZN => n1922);
   U2625 : OAI22_X1 port map( A1 => n8621, A2 => n8750, B1 => n8400, B2 => 
                           n8618, ZN => n1923);
   U2626 : OAI22_X1 port map( A1 => n8621, A2 => n8753, B1 => n8401, B2 => 
                           n3168, ZN => n1924);
   U2627 : OAI22_X1 port map( A1 => n8621, A2 => n8756, B1 => n8402, B2 => 
                           n3168, ZN => n1925);
   U2628 : OAI22_X1 port map( A1 => n8621, A2 => n8759, B1 => n8403, B2 => 
                           n3168, ZN => n1926);
   U2629 : OAI22_X1 port map( A1 => n8622, A2 => n8762, B1 => n8404, B2 => 
                           n8618, ZN => n1927);
   U2630 : OAI22_X1 port map( A1 => n8622, A2 => n8765, B1 => n8405, B2 => 
                           n8618, ZN => n1928);
   U2631 : OAI22_X1 port map( A1 => n8622, A2 => n8768, B1 => n8406, B2 => 
                           n8618, ZN => n1929);
   U2632 : OAI22_X1 port map( A1 => n8622, A2 => n8771, B1 => n8407, B2 => 
                           n8618, ZN => n1930);
   U2633 : OAI22_X1 port map( A1 => n8622, A2 => n8774, B1 => n8408, B2 => 
                           n8618, ZN => n1931);
   U2634 : OAI22_X1 port map( A1 => n8623, A2 => n8777, B1 => n8409, B2 => 
                           n8618, ZN => n1932);
   U2635 : OAI22_X1 port map( A1 => n8623, A2 => n8780, B1 => n8410, B2 => 
                           n8618, ZN => n1933);
   U2636 : OAI22_X1 port map( A1 => n8623, A2 => n8783, B1 => n8411, B2 => 
                           n8618, ZN => n1934);
   U2637 : OAI22_X1 port map( A1 => n8623, A2 => n8786, B1 => n8412, B2 => 
                           n8618, ZN => n1935);
   U2638 : OAI22_X1 port map( A1 => n8637, A2 => n8717, B1 => n6899, B2 => 
                           n8636, ZN => n1976);
   U2639 : OAI22_X1 port map( A1 => n8637, A2 => n8720, B1 => n6900, B2 => 
                           n8636, ZN => n1977);
   U2640 : OAI22_X1 port map( A1 => n8637, A2 => n8723, B1 => n6901, B2 => 
                           n8636, ZN => n1978);
   U2641 : OAI22_X1 port map( A1 => n8637, A2 => n8726, B1 => n6902, B2 => 
                           n8636, ZN => n1979);
   U2642 : OAI22_X1 port map( A1 => n8637, A2 => n8729, B1 => n6903, B2 => 
                           n8636, ZN => n1980);
   U2643 : OAI22_X1 port map( A1 => n8638, A2 => n8732, B1 => n6904, B2 => 
                           n8636, ZN => n1981);
   U2644 : OAI22_X1 port map( A1 => n8638, A2 => n8735, B1 => n6905, B2 => 
                           n8636, ZN => n1982);
   U2645 : OAI22_X1 port map( A1 => n8638, A2 => n8738, B1 => n6906, B2 => 
                           n8636, ZN => n1983);
   U2646 : OAI22_X1 port map( A1 => n8638, A2 => n8741, B1 => n6907, B2 => 
                           n8636, ZN => n1984);
   U2647 : OAI22_X1 port map( A1 => n8638, A2 => n8744, B1 => n6908, B2 => 
                           n8636, ZN => n1985);
   U2648 : OAI22_X1 port map( A1 => n8639, A2 => n8747, B1 => n6909, B2 => 
                           n8636, ZN => n1986);
   U2649 : OAI22_X1 port map( A1 => n8639, A2 => n8750, B1 => n6910, B2 => 
                           n8636, ZN => n1987);
   U2650 : OAI22_X1 port map( A1 => n8639, A2 => n8753, B1 => n6911, B2 => 
                           n3166, ZN => n1988);
   U2651 : OAI22_X1 port map( A1 => n8639, A2 => n8756, B1 => n6912, B2 => 
                           n3166, ZN => n1989);
   U2652 : OAI22_X1 port map( A1 => n8639, A2 => n8759, B1 => n6913, B2 => 
                           n3166, ZN => n1990);
   U2653 : OAI22_X1 port map( A1 => n8640, A2 => n8762, B1 => n6914, B2 => 
                           n8636, ZN => n1991);
   U2654 : OAI22_X1 port map( A1 => n8640, A2 => n8765, B1 => n6915, B2 => 
                           n8636, ZN => n1992);
   U2655 : OAI22_X1 port map( A1 => n8640, A2 => n8768, B1 => n6916, B2 => 
                           n8636, ZN => n1993);
   U2656 : OAI22_X1 port map( A1 => n8640, A2 => n8771, B1 => n6917, B2 => 
                           n8636, ZN => n1994);
   U2657 : OAI22_X1 port map( A1 => n8640, A2 => n8774, B1 => n6918, B2 => 
                           n8636, ZN => n1995);
   U2658 : OAI22_X1 port map( A1 => n8641, A2 => n8777, B1 => n6919, B2 => 
                           n8636, ZN => n1996);
   U2659 : OAI22_X1 port map( A1 => n8641, A2 => n8780, B1 => n6920, B2 => 
                           n8636, ZN => n1997);
   U2660 : OAI22_X1 port map( A1 => n8641, A2 => n8783, B1 => n6921, B2 => 
                           n8636, ZN => n1998);
   U2661 : OAI22_X1 port map( A1 => n8641, A2 => n8786, B1 => n6922, B2 => 
                           n8636, ZN => n1999);
   U2662 : OAI22_X1 port map( A1 => n8682, A2 => n8717, B1 => n8413, B2 => 
                           n8681, ZN => n2136);
   U2663 : OAI22_X1 port map( A1 => n8682, A2 => n8720, B1 => n8414, B2 => 
                           n8681, ZN => n2137);
   U2664 : OAI22_X1 port map( A1 => n8682, A2 => n8723, B1 => n8415, B2 => 
                           n8681, ZN => n2138);
   U2665 : OAI22_X1 port map( A1 => n8682, A2 => n8726, B1 => n8416, B2 => 
                           n8681, ZN => n2139);
   U2666 : OAI22_X1 port map( A1 => n8682, A2 => n8729, B1 => n8417, B2 => 
                           n8681, ZN => n2140);
   U2667 : OAI22_X1 port map( A1 => n8683, A2 => n8732, B1 => n8418, B2 => 
                           n8681, ZN => n2141);
   U2668 : OAI22_X1 port map( A1 => n8683, A2 => n8735, B1 => n8419, B2 => 
                           n8681, ZN => n2142);
   U2669 : OAI22_X1 port map( A1 => n8683, A2 => n8738, B1 => n8420, B2 => 
                           n8681, ZN => n2143);
   U2670 : OAI22_X1 port map( A1 => n8683, A2 => n8741, B1 => n8421, B2 => 
                           n8681, ZN => n2144);
   U2671 : OAI22_X1 port map( A1 => n8683, A2 => n8744, B1 => n8422, B2 => 
                           n8681, ZN => n2145);
   U2672 : OAI22_X1 port map( A1 => n8684, A2 => n8747, B1 => n8423, B2 => 
                           n8681, ZN => n2146);
   U2673 : OAI22_X1 port map( A1 => n8684, A2 => n8750, B1 => n8424, B2 => 
                           n8681, ZN => n2147);
   U2674 : OAI22_X1 port map( A1 => n8684, A2 => n8753, B1 => n8425, B2 => 
                           n3156, ZN => n2148);
   U2675 : OAI22_X1 port map( A1 => n8684, A2 => n8756, B1 => n8426, B2 => 
                           n3156, ZN => n2149);
   U2676 : OAI22_X1 port map( A1 => n8684, A2 => n8759, B1 => n8427, B2 => 
                           n3156, ZN => n2150);
   U2677 : OAI22_X1 port map( A1 => n8685, A2 => n8762, B1 => n8428, B2 => 
                           n8681, ZN => n2151);
   U2678 : OAI22_X1 port map( A1 => n8685, A2 => n8765, B1 => n8429, B2 => 
                           n8681, ZN => n2152);
   U2679 : OAI22_X1 port map( A1 => n8685, A2 => n8768, B1 => n8430, B2 => 
                           n8681, ZN => n2153);
   U2680 : OAI22_X1 port map( A1 => n8685, A2 => n8771, B1 => n8431, B2 => 
                           n8681, ZN => n2154);
   U2681 : OAI22_X1 port map( A1 => n8685, A2 => n8774, B1 => n8432, B2 => 
                           n8681, ZN => n2155);
   U2682 : OAI22_X1 port map( A1 => n8686, A2 => n8777, B1 => n8433, B2 => 
                           n8681, ZN => n2156);
   U2683 : OAI22_X1 port map( A1 => n8686, A2 => n8780, B1 => n8434, B2 => 
                           n8681, ZN => n2157);
   U2684 : OAI22_X1 port map( A1 => n8686, A2 => n8783, B1 => n8435, B2 => 
                           n8681, ZN => n2158);
   U2685 : OAI22_X1 port map( A1 => n8686, A2 => n8786, B1 => n8436, B2 => 
                           n8681, ZN => n2159);
   U2686 : NAND4_X1 port map( A1 => n2494, A2 => n2495, A3 => n2496, A4 => 
                           n2497, ZN => n3227);
   U2687 : AOI221_X1 port map( B1 => n8833, B2 => n3791, C1 => n8830, C2 => 
                           n3447, A => n2542, ZN => n2494);
   U2688 : AOI221_X1 port map( B1 => n8845, B2 => n6635, C1 => n8842, C2 => 
                           n6347, A => n2537, ZN => n2495);
   U2689 : NOR4_X1 port map( A1 => n2522, A2 => n2523, A3 => n2524, A4 => n2525
                           , ZN => n2496);
   U2690 : NAND4_X1 port map( A1 => n2545, A2 => n2546, A3 => n2547, A4 => 
                           n2548, ZN => n3226);
   U2691 : AOI221_X1 port map( B1 => n8833, B2 => n3792, C1 => n8830, C2 => 
                           n3448, A => n2562, ZN => n2545);
   U2692 : AOI221_X1 port map( B1 => n8845, B2 => n6636, C1 => n8842, C2 => 
                           n6348, A => n2561, ZN => n2546);
   U2693 : NOR4_X1 port map( A1 => n2557, A2 => n2558, A3 => n2559, A4 => n2560
                           , ZN => n2547);
   U2694 : NAND4_X1 port map( A1 => n2563, A2 => n2564, A3 => n2565, A4 => 
                           n2566, ZN => n3225);
   U2695 : AOI221_X1 port map( B1 => n8833, B2 => n3793, C1 => n8830, C2 => 
                           n3449, A => n2580, ZN => n2563);
   U2696 : AOI221_X1 port map( B1 => n8845, B2 => n6637, C1 => n8842, C2 => 
                           n6349, A => n2579, ZN => n2564);
   U2697 : NOR4_X1 port map( A1 => n2575, A2 => n2576, A3 => n2577, A4 => n2578
                           , ZN => n2565);
   U2698 : NAND4_X1 port map( A1 => n2581, A2 => n2582, A3 => n2583, A4 => 
                           n2584, ZN => n3224);
   U2699 : AOI221_X1 port map( B1 => n8833, B2 => n3794, C1 => n8830, C2 => 
                           n3450, A => n2598, ZN => n2581);
   U2700 : AOI221_X1 port map( B1 => n8845, B2 => n6638, C1 => n8842, C2 => 
                           n6350, A => n2597, ZN => n2582);
   U2701 : NOR4_X1 port map( A1 => n2593, A2 => n2594, A3 => n2595, A4 => n2596
                           , ZN => n2583);
   U2702 : NAND4_X1 port map( A1 => n2599, A2 => n2600, A3 => n2601, A4 => 
                           n2602, ZN => n3223);
   U2703 : AOI221_X1 port map( B1 => n8833, B2 => n3795, C1 => n8830, C2 => 
                           n3451, A => n2616, ZN => n2599);
   U2704 : AOI221_X1 port map( B1 => n8845, B2 => n6639, C1 => n8842, C2 => 
                           n6351, A => n2615, ZN => n2600);
   U2705 : NOR4_X1 port map( A1 => n2611, A2 => n2612, A3 => n2613, A4 => n2614
                           , ZN => n2601);
   U2706 : NAND4_X1 port map( A1 => n2617, A2 => n2618, A3 => n2619, A4 => 
                           n2620, ZN => n3222);
   U2707 : AOI221_X1 port map( B1 => n8833, B2 => n3796, C1 => n8830, C2 => 
                           n3452, A => n2634, ZN => n2617);
   U2708 : AOI221_X1 port map( B1 => n8845, B2 => n6640, C1 => n8842, C2 => 
                           n6352, A => n2633, ZN => n2618);
   U2709 : NOR4_X1 port map( A1 => n2629, A2 => n2630, A3 => n2631, A4 => n2632
                           , ZN => n2619);
   U2710 : NAND4_X1 port map( A1 => n2635, A2 => n2636, A3 => n2637, A4 => 
                           n2638, ZN => n3221);
   U2711 : AOI221_X1 port map( B1 => n8833, B2 => n3797, C1 => n8830, C2 => 
                           n3453, A => n2652, ZN => n2635);
   U2712 : AOI221_X1 port map( B1 => n8845, B2 => n6641, C1 => n8842, C2 => 
                           n6353, A => n2651, ZN => n2636);
   U2713 : NOR4_X1 port map( A1 => n2647, A2 => n2648, A3 => n2649, A4 => n2650
                           , ZN => n2637);
   U2714 : NAND4_X1 port map( A1 => n2653, A2 => n2654, A3 => n2655, A4 => 
                           n2656, ZN => n3220);
   U2715 : AOI221_X1 port map( B1 => n8833, B2 => n3798, C1 => n8830, C2 => 
                           n3454, A => n2670, ZN => n2653);
   U2716 : AOI221_X1 port map( B1 => n8845, B2 => n6642, C1 => n8842, C2 => 
                           n6354, A => n2669, ZN => n2654);
   U2717 : NOR4_X1 port map( A1 => n2665, A2 => n2666, A3 => n2667, A4 => n2668
                           , ZN => n2655);
   U2718 : NAND4_X1 port map( A1 => n2671, A2 => n2672, A3 => n2673, A4 => 
                           n2674, ZN => n3219);
   U2719 : AOI221_X1 port map( B1 => n8832, B2 => n3799, C1 => n8829, C2 => 
                           n3455, A => n2688, ZN => n2671);
   U2720 : AOI221_X1 port map( B1 => n8844, B2 => n6643, C1 => n8841, C2 => 
                           n6355, A => n2687, ZN => n2672);
   U2721 : NOR4_X1 port map( A1 => n2683, A2 => n2684, A3 => n2685, A4 => n2686
                           , ZN => n2673);
   U2722 : NAND4_X1 port map( A1 => n2689, A2 => n2690, A3 => n2691, A4 => 
                           n2692, ZN => n3218);
   U2723 : AOI221_X1 port map( B1 => n8832, B2 => n3800, C1 => n8829, C2 => 
                           n3456, A => n2706, ZN => n2689);
   U2724 : AOI221_X1 port map( B1 => n8844, B2 => n6644, C1 => n8841, C2 => 
                           n6356, A => n2705, ZN => n2690);
   U2725 : NOR4_X1 port map( A1 => n2701, A2 => n2702, A3 => n2703, A4 => n2704
                           , ZN => n2691);
   U2726 : NAND4_X1 port map( A1 => n2707, A2 => n2708, A3 => n2709, A4 => 
                           n2710, ZN => n3217);
   U2727 : AOI221_X1 port map( B1 => n8832, B2 => n3801, C1 => n8829, C2 => 
                           n3457, A => n2724, ZN => n2707);
   U2728 : AOI221_X1 port map( B1 => n8844, B2 => n6645, C1 => n8841, C2 => 
                           n6357, A => n2723, ZN => n2708);
   U2729 : NOR4_X1 port map( A1 => n2719, A2 => n2720, A3 => n2721, A4 => n2722
                           , ZN => n2709);
   U2730 : NAND4_X1 port map( A1 => n2725, A2 => n2726, A3 => n2727, A4 => 
                           n2728, ZN => n3216);
   U2731 : AOI221_X1 port map( B1 => n8832, B2 => n3802, C1 => n8829, C2 => 
                           n3458, A => n2742, ZN => n2725);
   U2732 : AOI221_X1 port map( B1 => n8844, B2 => n6646, C1 => n8841, C2 => 
                           n6358, A => n2741, ZN => n2726);
   U2733 : NOR4_X1 port map( A1 => n2737, A2 => n2738, A3 => n2739, A4 => n2740
                           , ZN => n2727);
   U2734 : NAND4_X1 port map( A1 => n2743, A2 => n2744, A3 => n2745, A4 => 
                           n2746, ZN => n3215);
   U2735 : AOI221_X1 port map( B1 => n8832, B2 => n3803, C1 => n8829, C2 => 
                           n3459, A => n2760, ZN => n2743);
   U2736 : AOI221_X1 port map( B1 => n8844, B2 => n6647, C1 => n8841, C2 => 
                           n6359, A => n2759, ZN => n2744);
   U2737 : NOR4_X1 port map( A1 => n2755, A2 => n2756, A3 => n2757, A4 => n2758
                           , ZN => n2745);
   U2738 : NAND4_X1 port map( A1 => n2761, A2 => n2762, A3 => n2763, A4 => 
                           n2764, ZN => n3214);
   U2739 : AOI221_X1 port map( B1 => n8832, B2 => n3804, C1 => n8829, C2 => 
                           n3460, A => n2778, ZN => n2761);
   U2740 : AOI221_X1 port map( B1 => n8844, B2 => n6648, C1 => n8841, C2 => 
                           n6360, A => n2777, ZN => n2762);
   U2741 : NOR4_X1 port map( A1 => n2773, A2 => n2774, A3 => n2775, A4 => n2776
                           , ZN => n2763);
   U2742 : NAND4_X1 port map( A1 => n2779, A2 => n2780, A3 => n2781, A4 => 
                           n2782, ZN => n3213);
   U2743 : AOI221_X1 port map( B1 => n8832, B2 => n3805, C1 => n8829, C2 => 
                           n3461, A => n2796, ZN => n2779);
   U2744 : AOI221_X1 port map( B1 => n8844, B2 => n6649, C1 => n8841, C2 => 
                           n6361, A => n2795, ZN => n2780);
   U2745 : NOR4_X1 port map( A1 => n2791, A2 => n2792, A3 => n2793, A4 => n2794
                           , ZN => n2781);
   U2746 : NAND4_X1 port map( A1 => n2797, A2 => n2798, A3 => n2799, A4 => 
                           n2800, ZN => n3212);
   U2747 : AOI221_X1 port map( B1 => n8832, B2 => n3806, C1 => n8829, C2 => 
                           n3462, A => n2814, ZN => n2797);
   U2748 : AOI221_X1 port map( B1 => n8844, B2 => n6650, C1 => n8841, C2 => 
                           n6362, A => n2813, ZN => n2798);
   U2749 : NOR4_X1 port map( A1 => n2809, A2 => n2810, A3 => n2811, A4 => n2812
                           , ZN => n2799);
   U2750 : NAND4_X1 port map( A1 => n2815, A2 => n2816, A3 => n2817, A4 => 
                           n2818, ZN => n3211);
   U2751 : AOI221_X1 port map( B1 => n8832, B2 => n3807, C1 => n8829, C2 => 
                           n3463, A => n2832, ZN => n2815);
   U2752 : AOI221_X1 port map( B1 => n8844, B2 => n6651, C1 => n8841, C2 => 
                           n6363, A => n2831, ZN => n2816);
   U2753 : NOR4_X1 port map( A1 => n2827, A2 => n2828, A3 => n2829, A4 => n2830
                           , ZN => n2817);
   U2754 : NAND4_X1 port map( A1 => n2833, A2 => n2834, A3 => n2835, A4 => 
                           n2836, ZN => n3210);
   U2755 : AOI221_X1 port map( B1 => n8832, B2 => n3808, C1 => n8829, C2 => 
                           n3464, A => n2850, ZN => n2833);
   U2756 : AOI221_X1 port map( B1 => n8844, B2 => n6652, C1 => n8841, C2 => 
                           n6364, A => n2849, ZN => n2834);
   U2757 : NOR4_X1 port map( A1 => n2845, A2 => n2846, A3 => n2847, A4 => n2848
                           , ZN => n2835);
   U2758 : NAND4_X1 port map( A1 => n2851, A2 => n2852, A3 => n2853, A4 => 
                           n2854, ZN => n3209);
   U2759 : AOI221_X1 port map( B1 => n8832, B2 => n3809, C1 => n8829, C2 => 
                           n3465, A => n2868, ZN => n2851);
   U2760 : AOI221_X1 port map( B1 => n8844, B2 => n6653, C1 => n8841, C2 => 
                           n6365, A => n2867, ZN => n2852);
   U2761 : NOR4_X1 port map( A1 => n2863, A2 => n2864, A3 => n2865, A4 => n2866
                           , ZN => n2853);
   U2762 : NAND4_X1 port map( A1 => n2869, A2 => n2870, A3 => n2871, A4 => 
                           n2872, ZN => n3208);
   U2763 : AOI221_X1 port map( B1 => n8832, B2 => n3810, C1 => n8829, C2 => 
                           n3466, A => n2886, ZN => n2869);
   U2764 : AOI221_X1 port map( B1 => n8844, B2 => n6654, C1 => n8841, C2 => 
                           n6366, A => n2885, ZN => n2870);
   U2765 : NOR4_X1 port map( A1 => n2881, A2 => n2882, A3 => n2883, A4 => n2884
                           , ZN => n2871);
   U2766 : NAND4_X1 port map( A1 => n2887, A2 => n2888, A3 => n2889, A4 => 
                           n2890, ZN => n3207);
   U2767 : AOI221_X1 port map( B1 => n8831, B2 => n3811, C1 => n8828, C2 => 
                           n3467, A => n2904, ZN => n2887);
   U2768 : AOI221_X1 port map( B1 => n8843, B2 => n6655, C1 => n8840, C2 => 
                           n6367, A => n2903, ZN => n2888);
   U2769 : NOR4_X1 port map( A1 => n2899, A2 => n2900, A3 => n2901, A4 => n2902
                           , ZN => n2889);
   U2770 : NAND4_X1 port map( A1 => n2905, A2 => n2906, A3 => n2907, A4 => 
                           n2908, ZN => n3206);
   U2771 : AOI221_X1 port map( B1 => n8831, B2 => n3812, C1 => n8828, C2 => 
                           n3468, A => n2922, ZN => n2905);
   U2772 : AOI221_X1 port map( B1 => n8843, B2 => n6656, C1 => n8840, C2 => 
                           n6368, A => n2921, ZN => n2906);
   U2773 : NOR4_X1 port map( A1 => n2917, A2 => n2918, A3 => n2919, A4 => n2920
                           , ZN => n2907);
   U2774 : NAND4_X1 port map( A1 => n2923, A2 => n2924, A3 => n2925, A4 => 
                           n2926, ZN => n3205);
   U2775 : AOI221_X1 port map( B1 => n8831, B2 => n3813, C1 => n8828, C2 => 
                           n3469, A => n2940, ZN => n2923);
   U2776 : AOI221_X1 port map( B1 => n8843, B2 => n6657, C1 => n8840, C2 => 
                           n6369, A => n2939, ZN => n2924);
   U2777 : NOR4_X1 port map( A1 => n2935, A2 => n2936, A3 => n2937, A4 => n2938
                           , ZN => n2925);
   U2778 : NAND4_X1 port map( A1 => n2941, A2 => n2942, A3 => n2943, A4 => 
                           n2944, ZN => n3204);
   U2779 : AOI221_X1 port map( B1 => n8831, B2 => n3814, C1 => n8828, C2 => 
                           n3470, A => n2958, ZN => n2941);
   U2780 : AOI221_X1 port map( B1 => n8843, B2 => n6658, C1 => n8840, C2 => 
                           n6370, A => n2957, ZN => n2942);
   U2781 : NOR4_X1 port map( A1 => n2953, A2 => n2954, A3 => n2955, A4 => n2956
                           , ZN => n2943);
   U2782 : NAND4_X1 port map( A1 => n2959, A2 => n2960, A3 => n2961, A4 => 
                           n2962, ZN => n3203);
   U2783 : AOI221_X1 port map( B1 => n8831, B2 => n3599, C1 => n8828, C2 => 
                           n3471, A => n2976, ZN => n2959);
   U2784 : AOI221_X1 port map( B1 => n8843, B2 => n6659, C1 => n8840, C2 => 
                           n6371, A => n2975, ZN => n2960);
   U2785 : NOR4_X1 port map( A1 => n2971, A2 => n2972, A3 => n2973, A4 => n2974
                           , ZN => n2961);
   U2786 : NAND4_X1 port map( A1 => n2977, A2 => n2978, A3 => n2979, A4 => 
                           n2980, ZN => n3202);
   U2787 : AOI221_X1 port map( B1 => n8831, B2 => n3600, C1 => n8828, C2 => 
                           n3472, A => n2994, ZN => n2977);
   U2788 : AOI221_X1 port map( B1 => n8843, B2 => n6660, C1 => n8840, C2 => 
                           n6372, A => n2993, ZN => n2978);
   U2789 : NOR4_X1 port map( A1 => n2989, A2 => n2990, A3 => n2991, A4 => n2992
                           , ZN => n2979);
   U2790 : NAND4_X1 port map( A1 => n2995, A2 => n2996, A3 => n2997, A4 => 
                           n2998, ZN => n3201);
   U2791 : AOI221_X1 port map( B1 => n8831, B2 => n3601, C1 => n8828, C2 => 
                           n3473, A => n3012, ZN => n2995);
   U2792 : AOI221_X1 port map( B1 => n8843, B2 => n6661, C1 => n8840, C2 => 
                           n6373, A => n3011, ZN => n2996);
   U2793 : NOR4_X1 port map( A1 => n3007, A2 => n3008, A3 => n3009, A4 => n3010
                           , ZN => n2997);
   U2794 : NAND4_X1 port map( A1 => n3013, A2 => n3014, A3 => n3015, A4 => 
                           n3016, ZN => n3200);
   U2795 : AOI221_X1 port map( B1 => n8831, B2 => n3602, C1 => n8828, C2 => 
                           n3474, A => n3030, ZN => n3013);
   U2796 : AOI221_X1 port map( B1 => n8843, B2 => n6662, C1 => n8840, C2 => 
                           n6374, A => n3029, ZN => n3014);
   U2797 : NOR4_X1 port map( A1 => n3025, A2 => n3026, A3 => n3027, A4 => n3028
                           , ZN => n3015);
   U2798 : NAND4_X1 port map( A1 => n3031, A2 => n3032, A3 => n3033, A4 => 
                           n3034, ZN => n3199);
   U2799 : AOI221_X1 port map( B1 => n8831, B2 => n3603, C1 => n8828, C2 => 
                           n3475, A => n3048, ZN => n3031);
   U2800 : AOI221_X1 port map( B1 => n8843, B2 => n6663, C1 => n8840, C2 => 
                           n6375, A => n3047, ZN => n3032);
   U2801 : NOR4_X1 port map( A1 => n3043, A2 => n3044, A3 => n3045, A4 => n3046
                           , ZN => n3033);
   U2802 : NAND4_X1 port map( A1 => n3049, A2 => n3050, A3 => n3051, A4 => 
                           n3052, ZN => n3198);
   U2803 : AOI221_X1 port map( B1 => n8831, B2 => n3604, C1 => n8828, C2 => 
                           n3476, A => n3066, ZN => n3049);
   U2804 : AOI221_X1 port map( B1 => n8843, B2 => n6664, C1 => n8840, C2 => 
                           n6376, A => n3065, ZN => n3050);
   U2805 : NOR4_X1 port map( A1 => n3061, A2 => n3062, A3 => n3063, A4 => n3064
                           , ZN => n3051);
   U2806 : NAND4_X1 port map( A1 => n3067, A2 => n3068, A3 => n3069, A4 => 
                           n3070, ZN => n3197);
   U2807 : AOI221_X1 port map( B1 => n8831, B2 => n3605, C1 => n8828, C2 => 
                           n3477, A => n3084, ZN => n3067);
   U2808 : AOI221_X1 port map( B1 => n8843, B2 => n6665, C1 => n8840, C2 => 
                           n6377, A => n3083, ZN => n3068);
   U2809 : NOR4_X1 port map( A1 => n3079, A2 => n3080, A3 => n3081, A4 => n3082
                           , ZN => n3069);
   U2810 : NAND4_X1 port map( A1 => n3085, A2 => n3086, A3 => n3087, A4 => 
                           n3088, ZN => n3196);
   U2811 : AOI221_X1 port map( B1 => n8831, B2 => n3606, C1 => n8828, C2 => 
                           n3478, A => n3114, ZN => n3085);
   U2812 : AOI221_X1 port map( B1 => n8843, B2 => n6666, C1 => n8840, C2 => 
                           n6378, A => n3113, ZN => n3086);
   U2813 : NOR4_X1 port map( A1 => n3108, A2 => n3109, A3 => n3110, A4 => n3111
                           , ZN => n3087);
   U2814 : NAND2_X1 port map( A1 => n849, A2 => n850, ZN => n3259);
   U2815 : NOR4_X1 port map( A1 => n851, A2 => n852, A3 => n853, A4 => n854, ZN
                           => n850);
   U2816 : NOR4_X1 port map( A1 => n876, A2 => n877, A3 => n878, A4 => n879, ZN
                           => n849);
   U2817 : OAI221_X1 port map( B1 => n6899, B2 => n8995, C1 => n6707, C2 => 
                           n8992, A => n867, ZN => n852);
   U2818 : NAND2_X1 port map( A1 => n900, A2 => n901, ZN => n3258);
   U2819 : NOR4_X1 port map( A1 => n902, A2 => n903, A3 => n904, A4 => n905, ZN
                           => n901);
   U2820 : NOR4_X1 port map( A1 => n910, A2 => n911, A3 => n912, A4 => n913, ZN
                           => n900);
   U2821 : OAI221_X1 port map( B1 => n6900, B2 => n8995, C1 => n6708, C2 => 
                           n8992, A => n908, ZN => n903);
   U2822 : NAND2_X1 port map( A1 => n918, A2 => n919, ZN => n3257);
   U2823 : NOR4_X1 port map( A1 => n920, A2 => n921, A3 => n922, A4 => n923, ZN
                           => n919);
   U2824 : NOR4_X1 port map( A1 => n928, A2 => n929, A3 => n930, A4 => n931, ZN
                           => n918);
   U2825 : OAI221_X1 port map( B1 => n6901, B2 => n8995, C1 => n6709, C2 => 
                           n8992, A => n926, ZN => n921);
   U2826 : NAND2_X1 port map( A1 => n936, A2 => n937, ZN => n3256);
   U2827 : NOR4_X1 port map( A1 => n938, A2 => n939, A3 => n940, A4 => n941, ZN
                           => n937);
   U2828 : NOR4_X1 port map( A1 => n946, A2 => n947, A3 => n948, A4 => n949, ZN
                           => n936);
   U2829 : OAI221_X1 port map( B1 => n6902, B2 => n8995, C1 => n6710, C2 => 
                           n8992, A => n944, ZN => n939);
   U2830 : NAND2_X1 port map( A1 => n954, A2 => n955, ZN => n3255);
   U2831 : NOR4_X1 port map( A1 => n956, A2 => n957, A3 => n958, A4 => n959, ZN
                           => n955);
   U2832 : NOR4_X1 port map( A1 => n964, A2 => n965, A3 => n966, A4 => n967, ZN
                           => n954);
   U2833 : OAI221_X1 port map( B1 => n6903, B2 => n8995, C1 => n6711, C2 => 
                           n8992, A => n962, ZN => n957);
   U2834 : NAND2_X1 port map( A1 => n972, A2 => n973, ZN => n3254);
   U2835 : NOR4_X1 port map( A1 => n974, A2 => n975, A3 => n976, A4 => n977, ZN
                           => n973);
   U2836 : NOR4_X1 port map( A1 => n982, A2 => n983, A3 => n984, A4 => n985, ZN
                           => n972);
   U2837 : OAI221_X1 port map( B1 => n6904, B2 => n8995, C1 => n6712, C2 => 
                           n8992, A => n980, ZN => n975);
   U2838 : NAND2_X1 port map( A1 => n990, A2 => n991, ZN => n3253);
   U2839 : NOR4_X1 port map( A1 => n992, A2 => n993, A3 => n994, A4 => n995, ZN
                           => n991);
   U2840 : NOR4_X1 port map( A1 => n1000, A2 => n1001, A3 => n1002, A4 => n1003
                           , ZN => n990);
   U2841 : OAI221_X1 port map( B1 => n6905, B2 => n8995, C1 => n6713, C2 => 
                           n8992, A => n998, ZN => n993);
   U2842 : NAND2_X1 port map( A1 => n1008, A2 => n1009, ZN => n3252);
   U2843 : NOR4_X1 port map( A1 => n1010, A2 => n1011, A3 => n1012, A4 => n1013
                           , ZN => n1009);
   U2844 : NOR4_X1 port map( A1 => n1018, A2 => n1019, A3 => n1020, A4 => n1021
                           , ZN => n1008);
   U2845 : OAI221_X1 port map( B1 => n6906, B2 => n8995, C1 => n6714, C2 => 
                           n8992, A => n1016, ZN => n1011);
   U2846 : NAND2_X1 port map( A1 => n1026, A2 => n1027, ZN => n3251);
   U2847 : NOR4_X1 port map( A1 => n1028, A2 => n1029, A3 => n1030, A4 => n1031
                           , ZN => n1027);
   U2848 : NOR4_X1 port map( A1 => n1036, A2 => n1037, A3 => n1038, A4 => n1039
                           , ZN => n1026);
   U2849 : OAI221_X1 port map( B1 => n6907, B2 => n8994, C1 => n6715, C2 => 
                           n8991, A => n1034, ZN => n1029);
   U2850 : NAND2_X1 port map( A1 => n1044, A2 => n1045, ZN => n3250);
   U2851 : NOR4_X1 port map( A1 => n1046, A2 => n1047, A3 => n1048, A4 => n1049
                           , ZN => n1045);
   U2852 : NOR4_X1 port map( A1 => n1054, A2 => n1055, A3 => n1056, A4 => n1057
                           , ZN => n1044);
   U2853 : OAI221_X1 port map( B1 => n6908, B2 => n8994, C1 => n6716, C2 => 
                           n8991, A => n1052, ZN => n1047);
   U2854 : NAND2_X1 port map( A1 => n1062, A2 => n1063, ZN => n3249);
   U2855 : NOR4_X1 port map( A1 => n1064, A2 => n1065, A3 => n1066, A4 => n1067
                           , ZN => n1063);
   U2856 : NOR4_X1 port map( A1 => n1072, A2 => n1073, A3 => n1074, A4 => n1075
                           , ZN => n1062);
   U2857 : OAI221_X1 port map( B1 => n6909, B2 => n8994, C1 => n6717, C2 => 
                           n8991, A => n1070, ZN => n1065);
   U2858 : NAND2_X1 port map( A1 => n1080, A2 => n1081, ZN => n3248);
   U2859 : NOR4_X1 port map( A1 => n1082, A2 => n1083, A3 => n1084, A4 => n1085
                           , ZN => n1081);
   U2860 : NOR4_X1 port map( A1 => n1090, A2 => n1091, A3 => n1092, A4 => n1093
                           , ZN => n1080);
   U2861 : OAI221_X1 port map( B1 => n6910, B2 => n8994, C1 => n6718, C2 => 
                           n8991, A => n1088, ZN => n1083);
   U2862 : NAND2_X1 port map( A1 => n1098, A2 => n1099, ZN => n3247);
   U2863 : NOR4_X1 port map( A1 => n1100, A2 => n1101, A3 => n1102, A4 => n1103
                           , ZN => n1099);
   U2864 : NOR4_X1 port map( A1 => n1108, A2 => n1109, A3 => n1110, A4 => n1111
                           , ZN => n1098);
   U2865 : OAI221_X1 port map( B1 => n6911, B2 => n8994, C1 => n6719, C2 => 
                           n8991, A => n1106, ZN => n1101);
   U2866 : NAND2_X1 port map( A1 => n1116, A2 => n1117, ZN => n3246);
   U2867 : NOR4_X1 port map( A1 => n1118, A2 => n1119, A3 => n1120, A4 => n1121
                           , ZN => n1117);
   U2868 : NOR4_X1 port map( A1 => n1126, A2 => n1127, A3 => n1128, A4 => n1129
                           , ZN => n1116);
   U2869 : OAI221_X1 port map( B1 => n6912, B2 => n8994, C1 => n6720, C2 => 
                           n8991, A => n1124, ZN => n1119);
   U2870 : NAND2_X1 port map( A1 => n1134, A2 => n1135, ZN => n3245);
   U2871 : NOR4_X1 port map( A1 => n1136, A2 => n1137, A3 => n1138, A4 => n1139
                           , ZN => n1135);
   U2872 : NOR4_X1 port map( A1 => n1144, A2 => n1145, A3 => n1146, A4 => n1147
                           , ZN => n1134);
   U2873 : OAI221_X1 port map( B1 => n6913, B2 => n8994, C1 => n6721, C2 => 
                           n8991, A => n1142, ZN => n1137);
   U2874 : NAND2_X1 port map( A1 => n1152, A2 => n1153, ZN => n3244);
   U2875 : NOR4_X1 port map( A1 => n1154, A2 => n1155, A3 => n1156, A4 => n1157
                           , ZN => n1153);
   U2876 : NOR4_X1 port map( A1 => n1162, A2 => n1163, A3 => n1164, A4 => n1165
                           , ZN => n1152);
   U2877 : OAI221_X1 port map( B1 => n6914, B2 => n8994, C1 => n6722, C2 => 
                           n8991, A => n1160, ZN => n1155);
   U2878 : NAND2_X1 port map( A1 => n1170, A2 => n1171, ZN => n3243);
   U2879 : NOR4_X1 port map( A1 => n1172, A2 => n1173, A3 => n1174, A4 => n1175
                           , ZN => n1171);
   U2880 : NOR4_X1 port map( A1 => n1180, A2 => n1181, A3 => n1182, A4 => n1183
                           , ZN => n1170);
   U2881 : OAI221_X1 port map( B1 => n6915, B2 => n8994, C1 => n6723, C2 => 
                           n8991, A => n1178, ZN => n1173);
   U2882 : NAND2_X1 port map( A1 => n1188, A2 => n1189, ZN => n3242);
   U2883 : NOR4_X1 port map( A1 => n1190, A2 => n1191, A3 => n1192, A4 => n1193
                           , ZN => n1189);
   U2884 : NOR4_X1 port map( A1 => n1198, A2 => n1199, A3 => n1200, A4 => n1201
                           , ZN => n1188);
   U2885 : OAI221_X1 port map( B1 => n6916, B2 => n8994, C1 => n6724, C2 => 
                           n8991, A => n1196, ZN => n1191);
   U2886 : NAND2_X1 port map( A1 => n1206, A2 => n1207, ZN => n3241);
   U2887 : NOR4_X1 port map( A1 => n1208, A2 => n1209, A3 => n1210, A4 => n1211
                           , ZN => n1207);
   U2888 : NOR4_X1 port map( A1 => n1216, A2 => n1217, A3 => n1218, A4 => n1219
                           , ZN => n1206);
   U2889 : OAI221_X1 port map( B1 => n6917, B2 => n8994, C1 => n6725, C2 => 
                           n8991, A => n1214, ZN => n1209);
   U2890 : NAND2_X1 port map( A1 => n1224, A2 => n1225, ZN => n3240);
   U2891 : NOR4_X1 port map( A1 => n1226, A2 => n1227, A3 => n1228, A4 => n1229
                           , ZN => n1225);
   U2892 : NOR4_X1 port map( A1 => n1234, A2 => n1235, A3 => n1236, A4 => n1237
                           , ZN => n1224);
   U2893 : OAI221_X1 port map( B1 => n6918, B2 => n8994, C1 => n6726, C2 => 
                           n8991, A => n1232, ZN => n1227);
   U2894 : NAND2_X1 port map( A1 => n1242, A2 => n1243, ZN => n3239);
   U2895 : NOR4_X1 port map( A1 => n1244, A2 => n1245, A3 => n1246, A4 => n1247
                           , ZN => n1243);
   U2896 : NOR4_X1 port map( A1 => n1252, A2 => n1253, A3 => n1254, A4 => n1255
                           , ZN => n1242);
   U2897 : OAI221_X1 port map( B1 => n6919, B2 => n8993, C1 => n6727, C2 => 
                           n8990, A => n1250, ZN => n1245);
   U2898 : NAND2_X1 port map( A1 => n1260, A2 => n1261, ZN => n3238);
   U2899 : NOR4_X1 port map( A1 => n1262, A2 => n1263, A3 => n1264, A4 => n1265
                           , ZN => n1261);
   U2900 : NOR4_X1 port map( A1 => n1270, A2 => n1271, A3 => n2296, A4 => n2297
                           , ZN => n1260);
   U2901 : OAI221_X1 port map( B1 => n6920, B2 => n8993, C1 => n6728, C2 => 
                           n8990, A => n1268, ZN => n1263);
   U2902 : NAND2_X1 port map( A1 => n2302, A2 => n2303, ZN => n3237);
   U2903 : NOR4_X1 port map( A1 => n2304, A2 => n2305, A3 => n2306, A4 => n2307
                           , ZN => n2303);
   U2904 : NOR4_X1 port map( A1 => n2312, A2 => n2313, A3 => n2314, A4 => n2315
                           , ZN => n2302);
   U2905 : OAI221_X1 port map( B1 => n6921, B2 => n8993, C1 => n6729, C2 => 
                           n8990, A => n2310, ZN => n2305);
   U2906 : NAND2_X1 port map( A1 => n2320, A2 => n2321, ZN => n3236);
   U2907 : NOR4_X1 port map( A1 => n2322, A2 => n2323, A3 => n2324, A4 => n2325
                           , ZN => n2321);
   U2908 : NOR4_X1 port map( A1 => n2330, A2 => n2331, A3 => n2332, A4 => n2333
                           , ZN => n2320);
   U2909 : OAI221_X1 port map( B1 => n6922, B2 => n8993, C1 => n6730, C2 => 
                           n8990, A => n2328, ZN => n2323);
   U2910 : NAND2_X1 port map( A1 => n2338, A2 => n2339, ZN => n3235);
   U2911 : NOR4_X1 port map( A1 => n2340, A2 => n2341, A3 => n2342, A4 => n2343
                           , ZN => n2339);
   U2912 : NOR4_X1 port map( A1 => n2348, A2 => n2349, A3 => n2350, A4 => n2351
                           , ZN => n2338);
   U2913 : OAI221_X1 port map( B1 => n6867, B2 => n8993, C1 => n6675, C2 => 
                           n8990, A => n2346, ZN => n2341);
   U2914 : NAND2_X1 port map( A1 => n2356, A2 => n2357, ZN => n3234);
   U2915 : NOR4_X1 port map( A1 => n2358, A2 => n2359, A3 => n2360, A4 => n2361
                           , ZN => n2357);
   U2916 : NOR4_X1 port map( A1 => n2366, A2 => n2367, A3 => n2368, A4 => n2369
                           , ZN => n2356);
   U2917 : OAI221_X1 port map( B1 => n6868, B2 => n8993, C1 => n6676, C2 => 
                           n8990, A => n2364, ZN => n2359);
   U2918 : NAND2_X1 port map( A1 => n2374, A2 => n2375, ZN => n3233);
   U2919 : NOR4_X1 port map( A1 => n2376, A2 => n2377, A3 => n2378, A4 => n2379
                           , ZN => n2375);
   U2920 : NOR4_X1 port map( A1 => n2384, A2 => n2385, A3 => n2386, A4 => n2387
                           , ZN => n2374);
   U2921 : OAI221_X1 port map( B1 => n6869, B2 => n8993, C1 => n6677, C2 => 
                           n8990, A => n2382, ZN => n2377);
   U2922 : NAND2_X1 port map( A1 => n2392, A2 => n2393, ZN => n3232);
   U2923 : NOR4_X1 port map( A1 => n2394, A2 => n2395, A3 => n2396, A4 => n2397
                           , ZN => n2393);
   U2924 : NOR4_X1 port map( A1 => n2402, A2 => n2403, A3 => n2404, A4 => n2405
                           , ZN => n2392);
   U2925 : OAI221_X1 port map( B1 => n6870, B2 => n8993, C1 => n6678, C2 => 
                           n8990, A => n2400, ZN => n2395);
   U2926 : NAND2_X1 port map( A1 => n2410, A2 => n2411, ZN => n3231);
   U2927 : NOR4_X1 port map( A1 => n2412, A2 => n2413, A3 => n2414, A4 => n2415
                           , ZN => n2411);
   U2928 : NOR4_X1 port map( A1 => n2420, A2 => n2421, A3 => n2422, A4 => n2423
                           , ZN => n2410);
   U2929 : OAI221_X1 port map( B1 => n6871, B2 => n8993, C1 => n6679, C2 => 
                           n8990, A => n2418, ZN => n2413);
   U2930 : NAND2_X1 port map( A1 => n2428, A2 => n2429, ZN => n3230);
   U2931 : NOR4_X1 port map( A1 => n2430, A2 => n2431, A3 => n2432, A4 => n2433
                           , ZN => n2429);
   U2932 : NOR4_X1 port map( A1 => n2438, A2 => n2439, A3 => n2440, A4 => n2441
                           , ZN => n2428);
   U2933 : OAI221_X1 port map( B1 => n6872, B2 => n8993, C1 => n6680, C2 => 
                           n8990, A => n2436, ZN => n2431);
   U2934 : NAND2_X1 port map( A1 => n2446, A2 => n2447, ZN => n3229);
   U2935 : NOR4_X1 port map( A1 => n2448, A2 => n2449, A3 => n2450, A4 => n2451
                           , ZN => n2447);
   U2936 : NOR4_X1 port map( A1 => n2456, A2 => n2457, A3 => n2458, A4 => n2459
                           , ZN => n2446);
   U2937 : OAI221_X1 port map( B1 => n6873, B2 => n8993, C1 => n6681, C2 => 
                           n8990, A => n2454, ZN => n2449);
   U2938 : NAND2_X1 port map( A1 => n2464, A2 => n2465, ZN => n3228);
   U2939 : NOR4_X1 port map( A1 => n2466, A2 => n2467, A3 => n2468, A4 => n2469
                           , ZN => n2465);
   U2940 : NOR4_X1 port map( A1 => n2484, A2 => n2485, A3 => n2486, A4 => n2487
                           , ZN => n2464);
   U2941 : OAI221_X1 port map( B1 => n6874, B2 => n8993, C1 => n6682, C2 => 
                           n8990, A => n2481, ZN => n2467);
   U2942 : NOR3_X1 port map( A1 => n845, A2 => ADD_RD2(2), A3 => n844, ZN => 
                           n2474);
   U2943 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(2), ZN => n3112);
   U2944 : NAND4_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => WR, A4 =>
                           ENABLE, ZN => n3183);
   U2945 : NAND4_X1 port map( A1 => ADD_WR(4), A2 => WR, A3 => ENABLE, A4 => 
                           n835, ZN => n3174);
   U2946 : NAND4_X1 port map( A1 => ADD_WR(3), A2 => WR, A3 => ENABLE, A4 => 
                           n834, ZN => n3165);
   U2947 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(4), A3 => n840, ZN
                           => n3105);
   U2948 : NOR3_X1 port map( A1 => n840, A2 => ADD_RD1(2), A3 => n839, ZN => 
                           n3107);
   U2949 : NOR3_X1 port map( A1 => n839, A2 => ADD_RD1(3), A3 => n841, ZN => 
                           n3097);
   U2950 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(3), A3 => n839, ZN
                           => n3106);
   U2951 : NAND4_X1 port map( A1 => WR, A2 => ENABLE, A3 => n835, A4 => n834, 
                           ZN => n3148);
   U2952 : NOR3_X1 port map( A1 => n844, A2 => ADD_RD2(3), A3 => n846, ZN => 
                           n2479);
   U2953 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n846, ZN
                           => n2491);
   U2954 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n841, ZN
                           => n3100);
   U2955 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(2), ZN => n2476);
   U2956 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(4), A3 => n845, ZN
                           => n2482);
   U2957 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(3), A3 => n844, ZN
                           => n2478);
   U2958 : INV_X1 port map( A => RESET, ZN => n833);
   U2959 : INV_X1 port map( A => ADD_RD2(2), ZN => n846);
   U2960 : INV_X1 port map( A => ADD_RD1(2), ZN => n841);
   U2961 : INV_X1 port map( A => ADD_RD2(3), ZN => n845);
   U2962 : INV_X1 port map( A => ADD_RD1(3), ZN => n840);
   U2963 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n9021, ZN => n3140);
   U2964 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n9021, ZN => n3138);
   U2965 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n9021, ZN => n3137);
   U2966 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n9021, ZN => n3136);
   U2967 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n9021, ZN => n3135);
   U2968 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n9021, ZN => n3134);
   U2969 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n9021, ZN => n3133);
   U2970 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n9021, ZN => n3132);
   U2971 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n9021, ZN => n3131);
   U2972 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n9021, ZN => n3130);
   U2973 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n9021, ZN => n3129);
   U2974 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n9021, ZN => n3128);
   U2975 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n9020, ZN => n3127);
   U2976 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n9020, ZN => n3126);
   U2977 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n9020, ZN => n3125);
   U2978 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n9020, ZN => n3124);
   U2979 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n9020, ZN => n3123);
   U2980 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n9020, ZN => n3122);
   U2981 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n9020, ZN => n3121);
   U2982 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n9020, ZN => n3120);
   U2983 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n9020, ZN => n3119);
   U2984 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n9020, ZN => n3118);
   U2985 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n9020, ZN => n3117);
   U2986 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n9020, ZN => n3115);
   U2987 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n9022, ZN => n3147);
   U2988 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n9022, ZN => n3146);
   U2989 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n9022, ZN => n3145);
   U2990 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n9022, ZN => n3144);
   U2991 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n9022, ZN => n3143);
   U2992 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n9022, ZN => n3142);
   U2993 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n9022, ZN => n3141);
   U2994 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n9022, ZN => n3139);
   U2995 : INV_X1 port map( A => ADD_WR(2), ZN => n836);
   U2996 : INV_X1 port map( A => ADD_WR(0), ZN => n838);
   U2997 : INV_X1 port map( A => ADD_WR(1), ZN => n837);
   U2998 : INV_X1 port map( A => ADD_WR(3), ZN => n835);
   U2999 : INV_X1 port map( A => ADD_RD2(0), ZN => n848);
   U3000 : INV_X1 port map( A => ADD_RD1(0), ZN => n843);
   U3001 : INV_X1 port map( A => ADD_RD2(1), ZN => n847);
   U3002 : INV_X1 port map( A => ADD_RD1(1), ZN => n842);
   U3003 : CLKBUF_X1 port map( A => n833, Z => n9025);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4.all;

entity 
   address_converter_NBIT_WIDTH32_F3_M8_N8_depth80_address_width5_address_ext4 
   is

   port( address_port_read_one, address_port_read_two, address_port_write, 
         cwp_in : in std_logic_vector (3 downto 0);  address_port_read_one_out,
         address_port_read_two_out, address_port_write_out : out 
         std_logic_vector (4 downto 0));

end address_converter_NBIT_WIDTH32_F3_M8_N8_depth80_address_width5_address_ext4
   ;

architecture SYN_Behavioral of 
   address_converter_NBIT_WIDTH32_F3_M8_N8_depth80_address_width5_address_ext4 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal address_port_read_one_out_4_port, address_port_read_two_out_4_port, 
      address_port_write_out_4_port : std_logic;

begin
   address_port_read_one_out <= ( address_port_read_one_out_4_port, 
      address_port_read_one(3), address_port_read_one(2), 
      address_port_read_one(1), address_port_read_one(0) );
   address_port_read_two_out <= ( address_port_read_two_out_4_port, 
      address_port_read_two(3), address_port_read_two(2), 
      address_port_read_two(1), address_port_read_two(0) );
   address_port_write_out <= ( address_port_write_out_4_port, 
      address_port_write(3), address_port_write(2), address_port_write(1), 
      address_port_write(0) );
   
   U3 : AND2_X1 port map( A1 => address_port_read_two(3), A2 => cwp_in(0), ZN 
                           => address_port_read_two_out_4_port);
   U4 : AND2_X1 port map( A1 => address_port_read_one(3), A2 => cwp_in(0), ZN 
                           => address_port_read_one_out_4_port);
   U5 : AND2_X1 port map( A1 => cwp_in(0), A2 => address_port_write(3), ZN => 
                           address_port_write_out_4_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4.all;

entity 
   register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4 
   is

   port( data_in_port_w : in std_logic_vector (31 downto 0);  data_out_port_a, 
         data_out_port_b : out std_logic_vector (31 downto 0);  
         address_port_read_one, address_port_read_two, address_port_write : in 
         std_logic_vector (3 downto 0);  r_signal_port_a, r_signal_port_b, 
         w_signal, clock, reset, enable, call, ret, mmu_ack : in std_logic;  
         cwp_out, swp_out : out std_logic_vector (3 downto 0);  fill, spill : 
         out std_logic);

end register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4;

architecture SYN_struct of 
   register_file_windowed_width_word32_F_reg3_m8_n8_address_ext4_log_port_rf4 
   is

   component control_unit
      port( clock, reset, call, ret, mmu_ack : in std_logic;  cwp_out, swp_out 
            : out std_logic_vector (3 downto 0);  fill, spill : out std_logic);
   end component;
   
   component register_file_NBIT32_NADDRESS5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      address_converter_NBIT_WIDTH32_F3_M8_N8_depth80_address_width5_address_ext4
      port( address_port_read_one, address_port_read_two, address_port_write, 
            cwp_in : in std_logic_vector (3 downto 0);  
            address_port_read_one_out, address_port_read_two_out, 
            address_port_write_out : out std_logic_vector (4 downto 0));
   end component;
   
   signal cwp_out_3_port, cwp_out_2_port, cwp_out_1_port, cwp_out_0_port, 
      swp_out_1_port, swp_out_0_port, address_port_read_one_out_4_port, 
      address_port_read_one_out_3_port, address_port_read_one_out_2_port, 
      address_port_read_one_out_1_port, address_port_read_one_out_0_port, 
      address_port_read_two_out_4_port, address_port_read_two_out_3_port, 
      address_port_read_two_out_2_port, address_port_read_two_out_1_port, 
      address_port_read_two_out_0_port, address_port_write_out_4_port, 
      address_port_write_out_3_port, address_port_write_out_2_port, 
      address_port_write_out_1_port, address_port_write_out_0_port, 
      swp_out_2_port, n_1448, n_1449 : std_logic;

begin
   cwp_out <= ( cwp_out_3_port, cwp_out_2_port, cwp_out_1_port, cwp_out_0_port 
      );
   swp_out <= ( swp_out_2_port, swp_out_2_port, swp_out_1_port, swp_out_0_port 
      );
   
   AC : 
                           address_converter_NBIT_WIDTH32_F3_M8_N8_depth80_address_width5_address_ext4 
                           port map( address_port_read_one(3) => 
                           address_port_read_one(3), address_port_read_one(2) 
                           => address_port_read_one(2), 
                           address_port_read_one(1) => address_port_read_one(1)
                           , address_port_read_one(0) => 
                           address_port_read_one(0), address_port_read_two(3) 
                           => address_port_read_two(3), 
                           address_port_read_two(2) => address_port_read_two(2)
                           , address_port_read_two(1) => 
                           address_port_read_two(1), address_port_read_two(0) 
                           => address_port_read_two(0), address_port_write(3) 
                           => address_port_write(3), address_port_write(2) => 
                           address_port_write(2), address_port_write(1) => 
                           address_port_write(1), address_port_write(0) => 
                           address_port_write(0), cwp_in(3) => cwp_out_3_port, 
                           cwp_in(2) => cwp_out_2_port, cwp_in(1) => 
                           cwp_out_1_port, cwp_in(0) => cwp_out_0_port, 
                           address_port_read_one_out(4) => 
                           address_port_read_one_out_4_port, 
                           address_port_read_one_out(3) => 
                           address_port_read_one_out_3_port, 
                           address_port_read_one_out(2) => 
                           address_port_read_one_out_2_port, 
                           address_port_read_one_out(1) => 
                           address_port_read_one_out_1_port, 
                           address_port_read_one_out(0) => 
                           address_port_read_one_out_0_port, 
                           address_port_read_two_out(4) => 
                           address_port_read_two_out_4_port, 
                           address_port_read_two_out(3) => 
                           address_port_read_two_out_3_port, 
                           address_port_read_two_out(2) => 
                           address_port_read_two_out_2_port, 
                           address_port_read_two_out(1) => 
                           address_port_read_two_out_1_port, 
                           address_port_read_two_out(0) => 
                           address_port_read_two_out_0_port, 
                           address_port_write_out(4) => 
                           address_port_write_out_4_port, 
                           address_port_write_out(3) => 
                           address_port_write_out_3_port, 
                           address_port_write_out(2) => 
                           address_port_write_out_2_port, 
                           address_port_write_out(1) => 
                           address_port_write_out_1_port, 
                           address_port_write_out(0) => 
                           address_port_write_out_0_port);
   RF : register_file_NBIT32_NADDRESS5 port map( CLK => clock, RESET => reset, 
                           ENABLE => enable, RD1 => r_signal_port_a, RD2 => 
                           r_signal_port_b, WR => w_signal, ADD_WR(4) => 
                           address_port_write_out_4_port, ADD_WR(3) => 
                           address_port_write_out_3_port, ADD_WR(2) => 
                           address_port_write_out_2_port, ADD_WR(1) => 
                           address_port_write_out_1_port, ADD_WR(0) => 
                           address_port_write_out_0_port, ADD_RD1(4) => 
                           address_port_read_one_out_4_port, ADD_RD1(3) => 
                           address_port_read_one_out_3_port, ADD_RD1(2) => 
                           address_port_read_one_out_2_port, ADD_RD1(1) => 
                           address_port_read_one_out_1_port, ADD_RD1(0) => 
                           address_port_read_one_out_0_port, ADD_RD2(4) => 
                           address_port_read_two_out_4_port, ADD_RD2(3) => 
                           address_port_read_two_out_3_port, ADD_RD2(2) => 
                           address_port_read_two_out_2_port, ADD_RD2(1) => 
                           address_port_read_two_out_1_port, ADD_RD2(0) => 
                           address_port_read_two_out_0_port, DATAIN(31) => 
                           data_in_port_w(31), DATAIN(30) => data_in_port_w(30)
                           , DATAIN(29) => data_in_port_w(29), DATAIN(28) => 
                           data_in_port_w(28), DATAIN(27) => data_in_port_w(27)
                           , DATAIN(26) => data_in_port_w(26), DATAIN(25) => 
                           data_in_port_w(25), DATAIN(24) => data_in_port_w(24)
                           , DATAIN(23) => data_in_port_w(23), DATAIN(22) => 
                           data_in_port_w(22), DATAIN(21) => data_in_port_w(21)
                           , DATAIN(20) => data_in_port_w(20), DATAIN(19) => 
                           data_in_port_w(19), DATAIN(18) => data_in_port_w(18)
                           , DATAIN(17) => data_in_port_w(17), DATAIN(16) => 
                           data_in_port_w(16), DATAIN(15) => data_in_port_w(15)
                           , DATAIN(14) => data_in_port_w(14), DATAIN(13) => 
                           data_in_port_w(13), DATAIN(12) => data_in_port_w(12)
                           , DATAIN(11) => data_in_port_w(11), DATAIN(10) => 
                           data_in_port_w(10), DATAIN(9) => data_in_port_w(9), 
                           DATAIN(8) => data_in_port_w(8), DATAIN(7) => 
                           data_in_port_w(7), DATAIN(6) => data_in_port_w(6), 
                           DATAIN(5) => data_in_port_w(5), DATAIN(4) => 
                           data_in_port_w(4), DATAIN(3) => data_in_port_w(3), 
                           DATAIN(2) => data_in_port_w(2), DATAIN(1) => 
                           data_in_port_w(1), DATAIN(0) => data_in_port_w(0), 
                           OUT1(31) => data_out_port_a(31), OUT1(30) => 
                           data_out_port_a(30), OUT1(29) => data_out_port_a(29)
                           , OUT1(28) => data_out_port_a(28), OUT1(27) => 
                           data_out_port_a(27), OUT1(26) => data_out_port_a(26)
                           , OUT1(25) => data_out_port_a(25), OUT1(24) => 
                           data_out_port_a(24), OUT1(23) => data_out_port_a(23)
                           , OUT1(22) => data_out_port_a(22), OUT1(21) => 
                           data_out_port_a(21), OUT1(20) => data_out_port_a(20)
                           , OUT1(19) => data_out_port_a(19), OUT1(18) => 
                           data_out_port_a(18), OUT1(17) => data_out_port_a(17)
                           , OUT1(16) => data_out_port_a(16), OUT1(15) => 
                           data_out_port_a(15), OUT1(14) => data_out_port_a(14)
                           , OUT1(13) => data_out_port_a(13), OUT1(12) => 
                           data_out_port_a(12), OUT1(11) => data_out_port_a(11)
                           , OUT1(10) => data_out_port_a(10), OUT1(9) => 
                           data_out_port_a(9), OUT1(8) => data_out_port_a(8), 
                           OUT1(7) => data_out_port_a(7), OUT1(6) => 
                           data_out_port_a(6), OUT1(5) => data_out_port_a(5), 
                           OUT1(4) => data_out_port_a(4), OUT1(3) => 
                           data_out_port_a(3), OUT1(2) => data_out_port_a(2), 
                           OUT1(1) => data_out_port_a(1), OUT1(0) => 
                           data_out_port_a(0), OUT2(31) => data_out_port_b(31),
                           OUT2(30) => data_out_port_b(30), OUT2(29) => 
                           data_out_port_b(29), OUT2(28) => data_out_port_b(28)
                           , OUT2(27) => data_out_port_b(27), OUT2(26) => 
                           data_out_port_b(26), OUT2(25) => data_out_port_b(25)
                           , OUT2(24) => data_out_port_b(24), OUT2(23) => 
                           data_out_port_b(23), OUT2(22) => data_out_port_b(22)
                           , OUT2(21) => data_out_port_b(21), OUT2(20) => 
                           data_out_port_b(20), OUT2(19) => data_out_port_b(19)
                           , OUT2(18) => data_out_port_b(18), OUT2(17) => 
                           data_out_port_b(17), OUT2(16) => data_out_port_b(16)
                           , OUT2(15) => data_out_port_b(15), OUT2(14) => 
                           data_out_port_b(14), OUT2(13) => data_out_port_b(13)
                           , OUT2(12) => data_out_port_b(12), OUT2(11) => 
                           data_out_port_b(11), OUT2(10) => data_out_port_b(10)
                           , OUT2(9) => data_out_port_b(9), OUT2(8) => 
                           data_out_port_b(8), OUT2(7) => data_out_port_b(7), 
                           OUT2(6) => data_out_port_b(6), OUT2(5) => 
                           data_out_port_b(5), OUT2(4) => data_out_port_b(4), 
                           OUT2(3) => data_out_port_b(3), OUT2(2) => 
                           data_out_port_b(2), OUT2(1) => data_out_port_b(1), 
                           OUT2(0) => data_out_port_b(0));
   CU : control_unit port map( clock => clock, reset => reset, call => call, 
                           ret => ret, mmu_ack => mmu_ack, cwp_out(3) => 
                           cwp_out_3_port, cwp_out(2) => cwp_out_2_port, 
                           cwp_out(1) => cwp_out_1_port, cwp_out(0) => 
                           cwp_out_0_port, swp_out(3) => n_1448, swp_out(2) => 
                           n_1449, swp_out(1) => swp_out_1_port, swp_out(0) => 
                           swp_out_0_port, fill => fill, spill => spill);
   swp_out_2_port <= '0';

end SYN_struct;
