library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity G_BLOCK is 
	
	
end G_BLOCK;

architecture BEHAVIORAL of G_BLOCK is
begin


end architecture BEHAVIORAL;