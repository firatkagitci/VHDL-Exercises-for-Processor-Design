package CONSTANTS is
   constant NumBit : integer := 32;	
   constant N_bit_address : integer := 5;
end CONSTANTS;
