library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;



entity PG_BLOCK is 

end G_BLOCK;

architecture BEHAVIORAL of PG_BLOCK is
begin

end architecture BEHAVIORAL;