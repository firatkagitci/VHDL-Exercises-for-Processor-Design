
module FD_0 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_127 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_126 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_125 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_124 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_123 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_122 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_121 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_120 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_119 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_118 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_117 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_116 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_115 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_114 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_113 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_112 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_111 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_110 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_109 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_108 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_107 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_106 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_105 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_104 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_103 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_102 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_101 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_100 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_99 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_98 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_97 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_GENERIC_NBIT32_0 ( D, CLK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET;
  wire   n7, n8, n9;

  FD_0 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n9), .Q(Q[0]) );
  FD_127 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n7), .Q(Q[1]) );
  FD_126 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n9), .Q(Q[2]) );
  FD_125 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n9), .Q(Q[3]) );
  FD_124 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n7), .Q(Q[4]) );
  FD_123 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n7), .Q(Q[5]) );
  FD_122 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n7), .Q(Q[6]) );
  FD_121 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n7), .Q(Q[7]) );
  FD_120 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n7), .Q(Q[8]) );
  FD_119 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n7), .Q(Q[9]) );
  FD_118 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n7), .Q(Q[10]) );
  FD_117 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n7), .Q(Q[11]) );
  FD_116 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n7), .Q(Q[12]) );
  FD_115 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n7), .Q(Q[13]) );
  FD_114 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n7), .Q(Q[14]) );
  FD_113 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n8), .Q(Q[15]) );
  FD_112 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n8), .Q(Q[16]) );
  FD_111 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n8), .Q(Q[17]) );
  FD_110 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n8), .Q(Q[18]) );
  FD_109 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n8), .Q(Q[19]) );
  FD_108 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n8), .Q(Q[20]) );
  FD_107 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n8), .Q(Q[21]) );
  FD_106 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n8), .Q(Q[22]) );
  FD_105 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n8), .Q(Q[23]) );
  FD_104 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n8), .Q(Q[24]) );
  FD_103 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n8), .Q(Q[25]) );
  FD_102 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n8), .Q(Q[26]) );
  FD_101 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n9), .Q(Q[27]) );
  FD_100 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n9), .Q(Q[28]) );
  FD_99 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n9), .Q(Q[29]) );
  FD_98 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n9), .Q(Q[30]) );
  FD_97 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n9), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n7) );
  BUF_X1 U2 ( .A(RESET), .Z(n8) );
  BUF_X1 U3 ( .A(RESET), .Z(n9) );
endmodule


module FD_96 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_95 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_94 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_93 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_92 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_91 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_90 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_89 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_88 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_87 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_86 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_85 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_84 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_83 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_82 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_81 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_80 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_79 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_78 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_77 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_76 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_75 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_74 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_73 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_72 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_71 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_70 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_69 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_68 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_67 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_66 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_65 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_GENERIC_NBIT32_1 ( D, CLK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET;
  wire   n7, n8, n9;

  FD_96 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n7), .Q(Q[0]) );
  FD_95 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n7), .Q(Q[1]) );
  FD_94 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n7), .Q(Q[2]) );
  FD_93 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n7), .Q(Q[3]) );
  FD_92 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n7), .Q(Q[4]) );
  FD_91 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n7), .Q(Q[5]) );
  FD_90 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n7), .Q(Q[6]) );
  FD_89 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n7), .Q(Q[7]) );
  FD_88 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n7), .Q(Q[8]) );
  FD_87 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n7), .Q(Q[9]) );
  FD_86 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n7), .Q(Q[10]) );
  FD_85 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n7), .Q(Q[11]) );
  FD_84 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n8), .Q(Q[12]) );
  FD_83 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n8), .Q(Q[13]) );
  FD_82 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n8), .Q(Q[14]) );
  FD_81 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n8), .Q(Q[15]) );
  FD_80 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n8), .Q(Q[16]) );
  FD_79 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n8), .Q(Q[17]) );
  FD_78 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n8), .Q(Q[18]) );
  FD_77 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n8), .Q(Q[19]) );
  FD_76 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n8), .Q(Q[20]) );
  FD_75 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n8), .Q(Q[21]) );
  FD_74 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n8), .Q(Q[22]) );
  FD_73 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n8), .Q(Q[23]) );
  FD_72 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n9), .Q(Q[24]) );
  FD_71 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n9), .Q(Q[25]) );
  FD_70 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n9), .Q(Q[26]) );
  FD_69 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n9), .Q(Q[27]) );
  FD_68 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n9), .Q(Q[28]) );
  FD_67 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n9), .Q(Q[29]) );
  FD_66 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n9), .Q(Q[30]) );
  FD_65 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n9), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n7) );
  BUF_X1 U2 ( .A(RESET), .Z(n8) );
  BUF_X1 U3 ( .A(RESET), .Z(n9) );
endmodule


module complement_NBIT64_0_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n223, n224, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n225, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301;

  XOR2_X1 U115 ( .A(n205), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U117 ( .A(n228), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U118 ( .A(n230), .B(B[60]), .Z(DIFF[60]) );
  NAND3_X1 U119 ( .A1(n299), .A2(n300), .A3(n232), .ZN(n230) );
  XOR2_X1 U120 ( .A(n226), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U121 ( .A(n234), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U122 ( .A(n235), .B(B[56]), .Z(DIFF[56]) );
  NAND3_X1 U123 ( .A1(n297), .A2(n298), .A3(n237), .ZN(n235) );
  XOR2_X1 U124 ( .A(n238), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U125 ( .A(n239), .B(B[52]), .Z(DIFF[52]) );
  NAND3_X1 U126 ( .A1(n295), .A2(n296), .A3(n241), .ZN(n239) );
  XOR2_X1 U127 ( .A(n242), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U128 ( .A(n233), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U129 ( .A(n243), .B(B[48]), .Z(DIFF[48]) );
  NAND3_X1 U130 ( .A1(n293), .A2(n294), .A3(n245), .ZN(n243) );
  XOR2_X1 U131 ( .A(n246), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U132 ( .A(n247), .B(B[44]), .Z(DIFF[44]) );
  NAND3_X1 U133 ( .A1(n291), .A2(n292), .A3(n249), .ZN(n247) );
  XOR2_X1 U134 ( .A(n250), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U135 ( .A(n251), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U136 ( .A(n204), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U137 ( .A(n255), .B(B[38]), .Z(DIFF[38]) );
  NAND3_X1 U138 ( .A1(n225), .A2(n288), .A3(n256), .ZN(n255) );
  XOR2_X1 U139 ( .A(n257), .B(n287), .Z(DIFF[37]) );
  XOR2_X1 U140 ( .A(n258), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U141 ( .A(n260), .B(B[32]), .Z(DIFF[32]) );
  NAND3_X1 U142 ( .A1(n202), .A2(n221), .A3(n220), .ZN(n260) );
  XOR2_X1 U144 ( .A(n264), .B(B[28]), .Z(DIFF[28]) );
  NAND3_X1 U145 ( .A1(n218), .A2(n219), .A3(n267), .ZN(n264) );
  XOR2_X1 U146 ( .A(n268), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U147 ( .A(n269), .B(B[24]), .Z(DIFF[24]) );
  NAND3_X1 U148 ( .A1(n216), .A2(n217), .A3(n271), .ZN(n269) );
  XOR2_X1 U149 ( .A(n272), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U150 ( .A(n273), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U151 ( .A(B[1]), .B(DIFF[0]), .Z(DIFF[1]) );
  XOR2_X1 U152 ( .A(n276), .B(B[18]), .Z(DIFF[18]) );
  NAND3_X1 U153 ( .A1(n213), .A2(n214), .A3(n277), .ZN(n276) );
  XOR2_X1 U154 ( .A(n278), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U155 ( .A(n279), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U156 ( .A(n285), .B(B[10]), .Z(DIFF[10]) );
  NOR3_X2 U3 ( .A1(n224), .A2(B[12]), .A3(n282), .ZN(n281) );
  NOR2_X2 U4 ( .A1(n273), .A2(n197), .ZN(n271) );
  NOR2_X2 U5 ( .A1(n269), .A2(n196), .ZN(n267) );
  NOR2_X1 U6 ( .A1(n258), .A2(B[35]), .ZN(n256) );
  OR2_X1 U7 ( .A1(B[24]), .A2(B[25]), .ZN(n196) );
  OR2_X1 U8 ( .A1(B[20]), .A2(B[21]), .ZN(n197) );
  OR2_X1 U9 ( .A1(B[15]), .A2(B[14]), .ZN(n198) );
  OR2_X1 U10 ( .A1(B[33]), .A2(B[32]), .ZN(n199) );
  XNOR2_X1 U11 ( .A(n200), .B(B[7]), .ZN(DIFF[7]) );
  NOR3_X1 U12 ( .A1(B[5]), .A2(B[6]), .A3(n226), .ZN(n200) );
  CLKBUF_X1 U13 ( .A(n265), .Z(n201) );
  NOR3_X1 U14 ( .A1(B[28]), .A2(B[29]), .A3(n264), .ZN(n202) );
  NOR3_X1 U15 ( .A1(B[28]), .A2(B[29]), .A3(n264), .ZN(n262) );
  CLKBUF_X1 U16 ( .A(n223), .Z(n203) );
  CLKBUF_X1 U17 ( .A(n254), .Z(n204) );
  OR3_X2 U18 ( .A1(n233), .A2(B[4]), .A3(n286), .ZN(n224) );
  OR3_X1 U19 ( .A1(n233), .A2(B[4]), .A3(n286), .ZN(n205) );
  CLKBUF_X1 U20 ( .A(B[0]), .Z(DIFF[0]) );
  NOR2_X1 U21 ( .A1(n279), .A2(n198), .ZN(n207) );
  AND2_X1 U22 ( .A1(n281), .A2(n208), .ZN(n277) );
  NOR2_X1 U23 ( .A1(B[13]), .A2(n198), .ZN(n208) );
  XNOR2_X1 U24 ( .A(n263), .B(n221), .ZN(DIFF[31]) );
  OR4_X1 U25 ( .A1(B[10]), .A2(B[11]), .A3(B[8]), .A4(B[9]), .ZN(n282) );
  OR2_X2 U26 ( .A1(n254), .A2(B[3]), .ZN(n233) );
  NOR3_X1 U27 ( .A1(n282), .A2(B[12]), .A3(n205), .ZN(n209) );
  NOR2_X1 U28 ( .A1(n260), .A2(n199), .ZN(n259) );
  NAND2_X1 U29 ( .A1(n253), .A2(n290), .ZN(n251) );
  NAND2_X1 U30 ( .A1(n241), .A2(n295), .ZN(n242) );
  NAND2_X1 U31 ( .A1(n245), .A2(n293), .ZN(n246) );
  NAND2_X1 U32 ( .A1(n237), .A2(n297), .ZN(n238) );
  NAND2_X1 U33 ( .A1(n232), .A2(n299), .ZN(n234) );
  NAND2_X1 U34 ( .A1(n229), .A2(n301), .ZN(n228) );
  NAND2_X1 U35 ( .A1(n256), .A2(n225), .ZN(n257) );
  NOR3_X1 U36 ( .A1(B[44]), .A2(B[45]), .A3(n247), .ZN(n245) );
  NOR3_X1 U37 ( .A1(B[48]), .A2(B[49]), .A3(n243), .ZN(n241) );
  NOR3_X1 U38 ( .A1(B[52]), .A2(B[53]), .A3(n239), .ZN(n237) );
  NOR3_X1 U39 ( .A1(B[56]), .A2(B[57]), .A3(n235), .ZN(n232) );
  NOR3_X1 U40 ( .A1(B[60]), .A2(B[61]), .A3(n230), .ZN(n229) );
  NOR3_X1 U41 ( .A1(B[40]), .A2(B[41]), .A3(n251), .ZN(n249) );
  NOR2_X1 U42 ( .A1(n255), .A2(B[38]), .ZN(n253) );
  XNOR2_X1 U43 ( .A(B[53]), .B(n240), .ZN(DIFF[53]) );
  NOR2_X1 U44 ( .A1(B[52]), .A2(n239), .ZN(n240) );
  XNOR2_X1 U45 ( .A(B[36]), .B(n256), .ZN(DIFF[36]) );
  XNOR2_X1 U46 ( .A(B[41]), .B(n252), .ZN(DIFF[41]) );
  NOR2_X1 U47 ( .A1(B[40]), .A2(n251), .ZN(n252) );
  XNOR2_X1 U48 ( .A(B[54]), .B(n237), .ZN(DIFF[54]) );
  XNOR2_X1 U49 ( .A(n289), .B(n253), .ZN(DIFF[39]) );
  XNOR2_X1 U50 ( .A(B[57]), .B(n236), .ZN(DIFF[57]) );
  NOR2_X1 U51 ( .A1(B[56]), .A2(n235), .ZN(n236) );
  XNOR2_X1 U52 ( .A(B[58]), .B(n232), .ZN(DIFF[58]) );
  XNOR2_X1 U53 ( .A(B[61]), .B(n231), .ZN(DIFF[61]) );
  NOR2_X1 U54 ( .A1(B[60]), .A2(n230), .ZN(n231) );
  XNOR2_X1 U55 ( .A(B[62]), .B(n229), .ZN(DIFF[62]) );
  XNOR2_X1 U56 ( .A(B[33]), .B(n261), .ZN(DIFF[33]) );
  NOR2_X1 U57 ( .A1(B[32]), .A2(n260), .ZN(n261) );
  XNOR2_X1 U58 ( .A(B[49]), .B(n244), .ZN(DIFF[49]) );
  NOR2_X1 U59 ( .A1(B[48]), .A2(n243), .ZN(n244) );
  XNOR2_X1 U60 ( .A(B[45]), .B(n248), .ZN(DIFF[45]) );
  NOR2_X1 U61 ( .A1(B[44]), .A2(n247), .ZN(n248) );
  XNOR2_X1 U62 ( .A(B[50]), .B(n241), .ZN(DIFF[50]) );
  XNOR2_X1 U63 ( .A(B[46]), .B(n245), .ZN(DIFF[46]) );
  XNOR2_X1 U64 ( .A(B[21]), .B(n274), .ZN(DIFF[21]) );
  NOR2_X1 U65 ( .A1(B[20]), .A2(n273), .ZN(n274) );
  XNOR2_X1 U66 ( .A(B[19]), .B(n275), .ZN(DIFF[19]) );
  XNOR2_X1 U67 ( .A(B[15]), .B(n280), .ZN(DIFF[15]) );
  XNOR2_X1 U68 ( .A(B[12]), .B(n283), .ZN(DIFF[12]) );
  NOR2_X1 U69 ( .A1(n205), .A2(n282), .ZN(n283) );
  NOR2_X1 U70 ( .A1(n276), .A2(B[18]), .ZN(n275) );
  NOR2_X1 U71 ( .A1(B[14]), .A2(n279), .ZN(n280) );
  XNOR2_X1 U72 ( .A(B[6]), .B(n227), .ZN(DIFF[6]) );
  NOR2_X1 U73 ( .A1(B[5]), .A2(n226), .ZN(n227) );
  OR3_X1 U74 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n286) );
  NOR2_X1 U75 ( .A1(n224), .A2(B[8]), .ZN(n223) );
  XNOR2_X1 U76 ( .A(B[25]), .B(n270), .ZN(DIFF[25]) );
  XNOR2_X1 U77 ( .A(B[29]), .B(n266), .ZN(DIFF[29]) );
  NOR2_X1 U78 ( .A1(B[28]), .A2(n264), .ZN(n266) );
  OR2_X1 U79 ( .A1(n233), .A2(B[4]), .ZN(n226) );
  NAND2_X1 U80 ( .A1(n275), .A2(n215), .ZN(n273) );
  XNOR2_X1 U81 ( .A(B[13]), .B(n209), .ZN(DIFF[13]) );
  NAND2_X1 U82 ( .A1(n281), .A2(n212), .ZN(n279) );
  XNOR2_X1 U83 ( .A(B[42]), .B(n249), .ZN(DIFF[42]) );
  NAND2_X1 U84 ( .A1(n249), .A2(n291), .ZN(n250) );
  NOR2_X1 U85 ( .A1(B[24]), .A2(n269), .ZN(n270) );
  XNOR2_X1 U86 ( .A(B[22]), .B(n271), .ZN(DIFF[22]) );
  NAND2_X1 U87 ( .A1(n271), .A2(n216), .ZN(n272) );
  NOR2_X1 U88 ( .A1(B[10]), .A2(n285), .ZN(n284) );
  XNOR2_X1 U89 ( .A(n284), .B(B[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U90 ( .A(B[9]), .B(n203), .ZN(DIFF[9]) );
  NAND2_X1 U91 ( .A1(n223), .A2(n211), .ZN(n285) );
  XNOR2_X1 U92 ( .A(n201), .B(B[2]), .ZN(DIFF[2]) );
  NAND2_X1 U93 ( .A1(n265), .A2(n210), .ZN(n254) );
  XNOR2_X1 U94 ( .A(B[34]), .B(n259), .ZN(DIFF[34]) );
  NAND2_X1 U95 ( .A1(n259), .A2(n222), .ZN(n258) );
  XNOR2_X1 U96 ( .A(n202), .B(B[30]), .ZN(DIFF[30]) );
  NAND2_X1 U97 ( .A1(n262), .A2(n220), .ZN(n263) );
  XNOR2_X1 U98 ( .A(B[26]), .B(n267), .ZN(DIFF[26]) );
  NAND2_X1 U99 ( .A1(n267), .A2(n218), .ZN(n268) );
  NAND2_X1 U100 ( .A1(n207), .A2(n213), .ZN(n278) );
  XNOR2_X1 U101 ( .A(B[16]), .B(n207), .ZN(DIFF[16]) );
  NOR2_X1 U102 ( .A1(B[1]), .A2(B[0]), .ZN(n265) );
  INV_X1 U103 ( .A(B[2]), .ZN(n210) );
  INV_X1 U104 ( .A(B[9]), .ZN(n211) );
  INV_X1 U105 ( .A(B[13]), .ZN(n212) );
  INV_X1 U106 ( .A(B[16]), .ZN(n213) );
  INV_X1 U107 ( .A(B[17]), .ZN(n214) );
  INV_X1 U108 ( .A(B[19]), .ZN(n215) );
  INV_X1 U109 ( .A(B[22]), .ZN(n216) );
  INV_X1 U110 ( .A(B[23]), .ZN(n217) );
  INV_X1 U111 ( .A(B[26]), .ZN(n218) );
  INV_X1 U112 ( .A(B[27]), .ZN(n219) );
  INV_X1 U113 ( .A(B[30]), .ZN(n220) );
  INV_X1 U114 ( .A(B[31]), .ZN(n221) );
  INV_X1 U116 ( .A(B[34]), .ZN(n222) );
  INV_X1 U143 ( .A(B[36]), .ZN(n225) );
  INV_X1 U157 ( .A(n288), .ZN(n287) );
  INV_X1 U158 ( .A(B[37]), .ZN(n288) );
  INV_X1 U159 ( .A(n290), .ZN(n289) );
  INV_X1 U160 ( .A(B[39]), .ZN(n290) );
  INV_X1 U161 ( .A(B[42]), .ZN(n291) );
  INV_X1 U162 ( .A(B[43]), .ZN(n292) );
  INV_X1 U163 ( .A(B[46]), .ZN(n293) );
  INV_X1 U164 ( .A(B[47]), .ZN(n294) );
  INV_X1 U165 ( .A(B[50]), .ZN(n295) );
  INV_X1 U166 ( .A(B[51]), .ZN(n296) );
  INV_X1 U167 ( .A(B[54]), .ZN(n297) );
  INV_X1 U168 ( .A(B[55]), .ZN(n298) );
  INV_X1 U169 ( .A(B[58]), .ZN(n299) );
  INV_X1 U170 ( .A(B[59]), .ZN(n300) );
  INV_X1 U171 ( .A(B[62]), .ZN(n301) );
endmodule


module complement_NBIT64_0 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_0_DW01_sub_4 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_31_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , net515275, net515254, net515252, net515239, net515229,
         net515161, net515160, net515159, net515059, net514770, net535378,
         net536671, net536728, net535981, net535381, net538516, net515178,
         net515177, n1, n2, n3, n4, n5, n14, n18, n19, n20, n21, n23, n24, n25,
         n26, n27, n28, n30, n31, n32, n34, n35, n36, n38, n39, n40, n43, n45,
         n47, n48, n53, n55, n57, n58, n62, n64, n66, n67, n71, n73, n75, n76,
         n78, n79, n80, n85, n86, n87, n88, n90, n91, n96, n97, n105, n111,
         n113, n115, n116, n117, n118, n124, n126, n128, n129, n130, n135,
         n136, n137, n138, n139, n140, n146, n147, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U16 ( .A(n178), .B(net515178), .Z(DIFF[18]) );
  XOR2_X1 U20 ( .A(n177), .B(net535981), .Z(DIFF[17]) );
  XOR2_X1 U22 ( .A(n175), .B(net536671), .Z(DIFF[15]) );
  NAND3_X1 U36 ( .A1(n166), .A2(n164), .A3(n4), .ZN(net515275) );
  XOR2_X1 U46 ( .A(n176), .B(net535381), .Z(DIFF[16]) );
  XOR2_X1 U63 ( .A(n20), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U65 ( .A(n21), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U67 ( .A(net536728), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U116 ( .A(n192), .B(n115), .Z(DIFF[32]) );
  XOR2_X1 U117 ( .A(n2), .B(n193), .Z(DIFF[33]) );
  XOR2_X1 U118 ( .A(n197), .B(n230), .Z(DIFF[36]) );
  XOR2_X1 U119 ( .A(n195), .B(n124), .Z(DIFF[34]) );
  XOR2_X1 U120 ( .A(n113), .B(n198), .Z(DIFF[37]) );
  XOR2_X1 U121 ( .A(n91), .B(n202), .Z(DIFF[40]) );
  XOR2_X1 U122 ( .A(n23), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U123 ( .A(n205), .B(n97), .Z(DIFF[42]) );
  XOR2_X1 U129 ( .A(n73), .B(n212), .Z(DIFF[48]) );
  XOR2_X1 U135 ( .A(n207), .B(n90), .Z(DIFF[44]) );
  XOR2_X1 U136 ( .A(n88), .B(n208), .Z(DIFF[45]) );
  XOR2_X1 U137 ( .A(n210), .B(n87), .Z(DIFF[46]) );
  XOR2_X1 U138 ( .A(n213), .B(n231), .Z(DIFF[49]) );
  XOR2_X1 U139 ( .A(n25), .B(n214), .Z(DIFF[50]) );
  XOR2_X1 U140 ( .A(n217), .B(n232), .Z(DIFF[53]) );
  XOR2_X1 U141 ( .A(n26), .B(n218), .Z(DIFF[54]) );
  XOR2_X1 U147 ( .A(n43), .B(B[61]), .Z(DIFF[61]) );
  XOR2_X1 U157 ( .A(n27), .B(n222), .Z(DIFF[58]) );
  XOR2_X1 U158 ( .A(n221), .B(n233), .Z(DIFF[57]) );
  XOR2_X1 U159 ( .A(n45), .B(n224), .Z(DIFF[60]) );
  XOR2_X1 U160 ( .A(n40), .B(n225), .Z(DIFF[62]) );
  XOR2_X1 U161 ( .A(n64), .B(n216), .Z(DIFF[52]) );
  XOR2_X1 U162 ( .A(n55), .B(n220), .Z(DIFF[56]) );
  XOR2_X1 U175 ( .A(n19), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U176 ( .A(n180), .B(n229), .Z(DIFF[20]) );
  XOR2_X1 U177 ( .A(n190), .B(n137), .Z(DIFF[30]) );
  XOR2_X1 U180 ( .A(n164), .B(n5), .Z(DIFF[4]) );
  XOR2_X1 U181 ( .A(n181), .B(n30), .Z(DIFF[21]) );
  XOR2_X1 U188 ( .A(n182), .B(n153), .Z(DIFF[22]) );
  XOR2_X1 U189 ( .A(n184), .B(n28), .Z(DIFF[24]) );
  XOR2_X1 U190 ( .A(n186), .B(n147), .Z(DIFF[26]) );
  XOR2_X1 U191 ( .A(n189), .B(n138), .Z(DIFF[29]) );
  XOR2_X1 U213 ( .A(n188), .B(n140), .Z(DIFF[28]) );
  XOR2_X1 U217 ( .A(n185), .B(n32), .Z(DIFF[25]) );
  NAND3_X1 U244 ( .A1(n222), .A2(n223), .A3(n221), .ZN(n48) );
  NAND3_X1 U245 ( .A1(n218), .A2(n219), .A3(n217), .ZN(n58) );
  NAND3_X1 U246 ( .A1(n214), .A2(n215), .A3(n213), .ZN(n67) );
  NAND3_X1 U247 ( .A1(n237), .A2(n24), .A3(n78), .ZN(n76) );
  NAND3_X1 U252 ( .A1(n162), .A2(n238), .A3(n161), .ZN(n105) );
  NAND3_X1 U258 ( .A1(n236), .A2(n31), .A3(n128), .ZN(n126) );
  OR4_X1 U3 ( .A1(B[6]), .A2(B[5]), .A3(B[4]), .A4(B[7]), .ZN(net514770) );
  XOR2_X1 U4 ( .A(n158), .B(n165), .Z(DIFF[5]) );
  AND2_X1 U5 ( .A1(n5), .A2(n164), .ZN(n158) );
  XOR2_X1 U6 ( .A(n159), .B(B[63]), .Z(DIFF[63]) );
  NAND2_X1 U7 ( .A1(n40), .A2(n225), .ZN(n159) );
  XOR2_X1 U8 ( .A(B[9]), .B(n160), .Z(DIFF[9]) );
  NAND2_X1 U9 ( .A1(n34), .A2(n5), .ZN(n160) );
  NOR2_X1 U10 ( .A1(n113), .A2(n198), .ZN(n111) );
  NOR2_X1 U11 ( .A1(n91), .A2(n85), .ZN(n90) );
  NOR2_X1 U12 ( .A1(n23), .A2(B[41]), .ZN(n97) );
  NOR2_X1 U13 ( .A1(n88), .A2(n208), .ZN(n87) );
  OR2_X1 U14 ( .A1(n202), .A2(n91), .ZN(n23) );
  INV_X1 U15 ( .A(n66), .ZN(n231) );
  INV_X1 U17 ( .A(n57), .ZN(n232) );
  INV_X1 U18 ( .A(n47), .ZN(n233) );
  NAND4_X1 U19 ( .A1(n203), .A2(n206), .A3(n205), .A4(n204), .ZN(n85) );
  NOR2_X1 U21 ( .A1(n2), .A2(n193), .ZN(n124) );
  NOR2_X1 U23 ( .A1(n75), .A2(n76), .ZN(n73) );
  NOR2_X1 U24 ( .A1(n79), .A2(n80), .ZN(n78) );
  INV_X1 U25 ( .A(n85), .ZN(n237) );
  NAND2_X1 U26 ( .A1(n24), .A2(n230), .ZN(n91) );
  INV_X1 U27 ( .A(n75), .ZN(n230) );
  NAND2_X1 U28 ( .A1(n73), .A2(n212), .ZN(n66) );
  NAND2_X1 U29 ( .A1(n230), .A2(n197), .ZN(n113) );
  NAND2_X1 U30 ( .A1(n207), .A2(n90), .ZN(n88) );
  AND2_X1 U31 ( .A1(n213), .A2(n231), .ZN(n25) );
  NOR2_X1 U32 ( .A1(n66), .A2(n67), .ZN(n64) );
  NOR2_X1 U33 ( .A1(n57), .A2(n58), .ZN(n55) );
  NOR2_X1 U34 ( .A1(n47), .A2(n48), .ZN(n45) );
  NAND2_X1 U35 ( .A1(n64), .A2(n216), .ZN(n57) );
  NAND2_X1 U37 ( .A1(n55), .A2(n220), .ZN(n47) );
  NAND2_X1 U38 ( .A1(n45), .A2(n224), .ZN(n43) );
  AND2_X1 U39 ( .A1(n217), .A2(n232), .ZN(n26) );
  AND2_X1 U40 ( .A1(n221), .A2(n233), .ZN(n27) );
  NAND2_X1 U41 ( .A1(n210), .A2(n211), .ZN(n79) );
  NAND2_X1 U42 ( .A1(n207), .A2(n209), .ZN(n80) );
  NAND2_X1 U43 ( .A1(n115), .A2(n116), .ZN(n75) );
  NOR2_X1 U44 ( .A1(n117), .A2(n118), .ZN(n116) );
  NAND2_X1 U45 ( .A1(n192), .A2(n196), .ZN(n117) );
  NAND2_X1 U47 ( .A1(n194), .A2(n195), .ZN(n118) );
  NAND2_X1 U48 ( .A1(n226), .A2(n166), .ZN(n36) );
  INV_X1 U49 ( .A(n38), .ZN(n226) );
  NAND2_X1 U50 ( .A1(n192), .A2(n115), .ZN(n2) );
  AND4_X1 U51 ( .A1(n197), .A2(n201), .A3(n200), .A4(n199), .ZN(n24) );
  NOR2_X1 U52 ( .A1(B[61]), .A2(n43), .ZN(n40) );
  XNOR2_X1 U53 ( .A(n215), .B(n71), .ZN(DIFF[51]) );
  NAND2_X1 U54 ( .A1(n214), .A2(n25), .ZN(n71) );
  NOR2_X1 U55 ( .A1(net515059), .A2(n126), .ZN(n115) );
  NOR2_X1 U56 ( .A1(n129), .A2(n130), .ZN(n128) );
  INV_X1 U57 ( .A(n135), .ZN(n236) );
  NAND2_X1 U58 ( .A1(n200), .A2(n111), .ZN(n21) );
  XNOR2_X1 U59 ( .A(n219), .B(n62), .ZN(DIFF[55]) );
  NAND2_X1 U60 ( .A1(n218), .A2(n26), .ZN(n62) );
  XNOR2_X1 U61 ( .A(n223), .B(n53), .ZN(DIFF[59]) );
  NAND2_X1 U62 ( .A1(n222), .A2(n27), .ZN(n53) );
  XNOR2_X1 U64 ( .A(n111), .B(B[38]), .ZN(DIFF[38]) );
  NAND2_X1 U66 ( .A1(n195), .A2(n124), .ZN(n20) );
  XNOR2_X1 U68 ( .A(n206), .B(n96), .ZN(DIFF[43]) );
  NAND2_X1 U69 ( .A1(n205), .A2(n97), .ZN(n96) );
  XNOR2_X1 U70 ( .A(n211), .B(n86), .ZN(DIFF[47]) );
  NAND2_X1 U71 ( .A1(n210), .A2(n87), .ZN(n86) );
  NOR2_X1 U72 ( .A1(net514770), .A2(B[8]), .ZN(n34) );
  XNOR2_X1 U73 ( .A(n39), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U74 ( .A1(n234), .A2(n38), .ZN(n39) );
  NOR2_X1 U75 ( .A1(n228), .A2(n135), .ZN(n140) );
  INV_X1 U76 ( .A(n28), .ZN(n228) );
  NAND2_X1 U77 ( .A1(n164), .A2(n165), .ZN(n38) );
  AND2_X1 U78 ( .A1(n31), .A2(n229), .ZN(n28) );
  AND2_X1 U79 ( .A1(n32), .A2(n185), .ZN(n147) );
  AND2_X1 U80 ( .A1(n30), .A2(n181), .ZN(n153) );
  INV_X1 U81 ( .A(net515059), .ZN(n229) );
  INV_X1 U82 ( .A(net515229), .ZN(n227) );
  AND2_X1 U83 ( .A1(net535381), .A2(n176), .ZN(net535981) );
  AND2_X1 U84 ( .A1(n229), .A2(n180), .ZN(n30) );
  XOR2_X1 U85 ( .A(n171), .B(net515252), .Z(DIFF[11]) );
  XNOR2_X1 U86 ( .A(n136), .B(n191), .ZN(DIFF[31]) );
  NAND2_X1 U87 ( .A1(n137), .A2(n190), .ZN(n136) );
  XNOR2_X1 U88 ( .A(n187), .B(n146), .ZN(DIFF[27]) );
  NAND2_X1 U89 ( .A1(n186), .A2(n147), .ZN(n146) );
  XNOR2_X1 U90 ( .A(n183), .B(n152), .ZN(DIFF[23]) );
  NAND2_X1 U91 ( .A1(n182), .A2(n153), .ZN(n152) );
  XNOR2_X1 U92 ( .A(n162), .B(n139), .ZN(DIFF[2]) );
  XNOR2_X1 U93 ( .A(n179), .B(net515177), .ZN(DIFF[19]) );
  NAND2_X1 U94 ( .A1(n178), .A2(net515178), .ZN(net515177) );
  AND3_X1 U95 ( .A1(n154), .A2(n227), .A3(n174), .ZN(net536671) );
  NAND4_X1 U96 ( .A1(n184), .A2(n187), .A3(n186), .A4(n185), .ZN(n135) );
  NOR2_X1 U97 ( .A1(B[13]), .A2(B[12]), .ZN(n154) );
  NAND2_X1 U98 ( .A1(net515239), .A2(n5), .ZN(net515229) );
  NOR2_X1 U99 ( .A1(n235), .A2(net514770), .ZN(net515239) );
  INV_X1 U100 ( .A(n1), .ZN(n235) );
  NOR2_X1 U101 ( .A1(n156), .A2(net515254), .ZN(net515252) );
  NAND2_X1 U102 ( .A1(n170), .A2(n169), .ZN(net515254) );
  NAND2_X1 U103 ( .A1(n34), .A2(n5), .ZN(n156) );
  XNOR2_X1 U104 ( .A(n155), .B(B[13]), .ZN(DIFF[13]) );
  NOR2_X1 U105 ( .A1(net515229), .A2(B[12]), .ZN(n155) );
  AND3_X1 U106 ( .A1(n171), .A2(n14), .A3(n170), .ZN(n1) );
  NOR2_X1 U107 ( .A1(B[9]), .A2(B[8]), .ZN(n14) );
  NAND2_X1 U108 ( .A1(net535381), .A2(net515159), .ZN(net515059) );
  NOR2_X1 U109 ( .A1(net515160), .A2(net515161), .ZN(net515159) );
  NAND2_X1 U110 ( .A1(n176), .A2(n179), .ZN(net515160) );
  NAND2_X1 U111 ( .A1(n177), .A2(n178), .ZN(net515161) );
  AND4_X1 U112 ( .A1(net538516), .A2(n3), .A3(n1), .A4(n5), .ZN(net535381) );
  AND4_X1 U113 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n3) );
  AND4_X1 U114 ( .A1(n164), .A2(n165), .A3(n166), .A4(n167), .ZN(net538516) );
  AND2_X1 U115 ( .A1(net535981), .A2(n177), .ZN(net515178) );
  INV_X1 U124 ( .A(n5), .ZN(n234) );
  AND2_X1 U125 ( .A1(n138), .A2(n189), .ZN(n137) );
  NAND2_X1 U126 ( .A1(n188), .A2(n189), .ZN(n130) );
  NAND2_X1 U127 ( .A1(n190), .A2(n191), .ZN(n129) );
  AND2_X1 U128 ( .A1(n140), .A2(n188), .ZN(n138) );
  AND2_X1 U130 ( .A1(n28), .A2(n184), .ZN(n32) );
  AND4_X1 U131 ( .A1(n180), .A2(n183), .A3(n182), .A4(n181), .ZN(n31) );
  AND2_X1 U132 ( .A1(n18), .A2(n5), .ZN(net535378) );
  NOR2_X1 U133 ( .A1(net515275), .A2(n157), .ZN(n18) );
  NAND2_X1 U134 ( .A1(n168), .A2(n165), .ZN(n157) );
  AND2_X1 U142 ( .A1(n169), .A2(n167), .ZN(n4) );
  NAND2_X1 U143 ( .A1(n227), .A2(n154), .ZN(n19) );
  XNOR2_X1 U144 ( .A(n35), .B(B[7]), .ZN(DIFF[7]) );
  NOR2_X1 U145 ( .A1(n234), .A2(n36), .ZN(n35) );
  XNOR2_X1 U146 ( .A(n172), .B(net515229), .ZN(DIFF[12]) );
  NAND2_X1 U148 ( .A1(net538516), .A2(n5), .ZN(net536728) );
  AND4_X2 U149 ( .A1(n162), .A2(n238), .A3(n163), .A4(n161), .ZN(n5) );
  XOR2_X1 U150 ( .A(net535378), .B(n170), .Z(DIFF[10]) );
  XNOR2_X1 U151 ( .A(n163), .B(n105), .ZN(DIFF[3]) );
  NAND2_X1 U152 ( .A1(n161), .A2(n238), .ZN(n139) );
  XNOR2_X1 U153 ( .A(\B[0] ), .B(n161), .ZN(DIFF[1]) );
  INV_X1 U154 ( .A(\B[0] ), .ZN(n238) );
  INV_X1 U155 ( .A(B[1]), .ZN(n161) );
  INV_X1 U156 ( .A(B[2]), .ZN(n162) );
  INV_X1 U163 ( .A(B[3]), .ZN(n163) );
  INV_X1 U164 ( .A(B[4]), .ZN(n164) );
  INV_X1 U165 ( .A(B[5]), .ZN(n165) );
  INV_X1 U166 ( .A(B[6]), .ZN(n166) );
  INV_X1 U167 ( .A(B[7]), .ZN(n167) );
  INV_X1 U168 ( .A(B[8]), .ZN(n168) );
  INV_X1 U169 ( .A(B[9]), .ZN(n169) );
  INV_X1 U170 ( .A(B[10]), .ZN(n170) );
  INV_X1 U171 ( .A(B[11]), .ZN(n171) );
  INV_X1 U172 ( .A(B[12]), .ZN(n172) );
  INV_X1 U173 ( .A(B[13]), .ZN(n173) );
  INV_X1 U174 ( .A(B[14]), .ZN(n174) );
  INV_X1 U178 ( .A(B[15]), .ZN(n175) );
  INV_X1 U179 ( .A(B[16]), .ZN(n176) );
  INV_X1 U182 ( .A(B[17]), .ZN(n177) );
  INV_X1 U183 ( .A(B[18]), .ZN(n178) );
  INV_X1 U184 ( .A(B[19]), .ZN(n179) );
  INV_X1 U185 ( .A(B[20]), .ZN(n180) );
  INV_X1 U186 ( .A(B[21]), .ZN(n181) );
  INV_X1 U187 ( .A(B[22]), .ZN(n182) );
  INV_X1 U192 ( .A(B[23]), .ZN(n183) );
  INV_X1 U193 ( .A(B[24]), .ZN(n184) );
  INV_X1 U194 ( .A(B[25]), .ZN(n185) );
  INV_X1 U195 ( .A(B[26]), .ZN(n186) );
  INV_X1 U196 ( .A(B[27]), .ZN(n187) );
  INV_X1 U197 ( .A(B[28]), .ZN(n188) );
  INV_X1 U198 ( .A(B[29]), .ZN(n189) );
  INV_X1 U199 ( .A(B[30]), .ZN(n190) );
  INV_X1 U200 ( .A(B[31]), .ZN(n191) );
  INV_X1 U201 ( .A(B[32]), .ZN(n192) );
  INV_X1 U202 ( .A(n194), .ZN(n193) );
  INV_X1 U203 ( .A(B[33]), .ZN(n194) );
  INV_X1 U204 ( .A(B[34]), .ZN(n195) );
  INV_X1 U205 ( .A(B[35]), .ZN(n196) );
  INV_X1 U206 ( .A(B[36]), .ZN(n197) );
  INV_X1 U207 ( .A(n199), .ZN(n198) );
  INV_X1 U208 ( .A(B[37]), .ZN(n199) );
  INV_X1 U209 ( .A(B[38]), .ZN(n200) );
  INV_X1 U210 ( .A(B[39]), .ZN(n201) );
  INV_X1 U211 ( .A(n203), .ZN(n202) );
  INV_X1 U212 ( .A(B[40]), .ZN(n203) );
  INV_X1 U214 ( .A(B[41]), .ZN(n204) );
  INV_X1 U215 ( .A(B[42]), .ZN(n205) );
  INV_X1 U216 ( .A(B[43]), .ZN(n206) );
  INV_X1 U218 ( .A(B[44]), .ZN(n207) );
  INV_X1 U219 ( .A(n209), .ZN(n208) );
  INV_X1 U220 ( .A(B[45]), .ZN(n209) );
  INV_X1 U221 ( .A(B[46]), .ZN(n210) );
  INV_X1 U222 ( .A(B[47]), .ZN(n211) );
  INV_X1 U223 ( .A(B[48]), .ZN(n212) );
  INV_X1 U224 ( .A(B[49]), .ZN(n213) );
  INV_X1 U225 ( .A(B[50]), .ZN(n214) );
  INV_X1 U226 ( .A(B[51]), .ZN(n215) );
  INV_X1 U227 ( .A(B[52]), .ZN(n216) );
  INV_X1 U228 ( .A(B[53]), .ZN(n217) );
  INV_X1 U229 ( .A(B[54]), .ZN(n218) );
  INV_X1 U230 ( .A(B[55]), .ZN(n219) );
  INV_X1 U231 ( .A(B[56]), .ZN(n220) );
  INV_X1 U232 ( .A(B[57]), .ZN(n221) );
  INV_X1 U233 ( .A(B[58]), .ZN(n222) );
  INV_X1 U234 ( .A(B[59]), .ZN(n223) );
  INV_X1 U235 ( .A(B[60]), .ZN(n224) );
  INV_X1 U236 ( .A(B[62]), .ZN(n225) );
endmodule


module complement_NBIT64_31 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_31_DW01_sub_7 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_30_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n291, n292, n293, n294, n295, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n290, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U114 ( .A(B[9]), .B(n233), .Z(DIFF[9]) );
  XOR2_X1 U115 ( .A(n208), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U116 ( .A(n235), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U117 ( .A(n238), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U118 ( .A(n240), .B(B[60]), .Z(DIFF[60]) );
  NAND3_X1 U119 ( .A1(n308), .A2(n309), .A3(n242), .ZN(n240) );
  XOR2_X1 U120 ( .A(n237), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U121 ( .A(n244), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U122 ( .A(n245), .B(B[56]), .Z(DIFF[56]) );
  NAND3_X1 U123 ( .A1(n306), .A2(n307), .A3(n247), .ZN(n245) );
  XOR2_X1 U124 ( .A(n248), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U125 ( .A(n249), .B(B[52]), .Z(DIFF[52]) );
  NAND3_X1 U126 ( .A1(n304), .A2(n305), .A3(n251), .ZN(n249) );
  XOR2_X1 U127 ( .A(n252), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U128 ( .A(n253), .B(B[48]), .Z(DIFF[48]) );
  NAND3_X1 U129 ( .A1(n302), .A2(n303), .A3(n255), .ZN(n253) );
  XOR2_X1 U130 ( .A(n256), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U131 ( .A(n257), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U132 ( .A(n260), .B(B[42]), .Z(DIFF[42]) );
  NAND3_X1 U133 ( .A1(n299), .A2(n300), .A3(n261), .ZN(n260) );
  XOR2_X1 U134 ( .A(n262), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U135 ( .A(n264), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U136 ( .A(n263), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U137 ( .A(n266), .B(B[36]), .Z(DIFF[36]) );
  XOR2_X1 U138 ( .A(n269), .B(B[34]), .Z(DIFF[34]) );
  NAND3_X1 U139 ( .A1(n290), .A2(n296), .A3(n270), .ZN(n269) );
  XOR2_X1 U141 ( .A(n272), .B(B[30]), .Z(DIFF[30]) );
  NAND3_X1 U142 ( .A1(n231), .A2(n232), .A3(n274), .ZN(n272) );
  XOR2_X1 U144 ( .A(n277), .B(B[26]), .Z(DIFF[26]) );
  NAND3_X1 U145 ( .A1(n229), .A2(n230), .A3(n279), .ZN(n277) );
  XOR2_X1 U147 ( .A(n281), .B(B[22]), .Z(DIFF[22]) );
  NAND3_X1 U148 ( .A1(n227), .A2(n228), .A3(n283), .ZN(n281) );
  XOR2_X1 U150 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U151 ( .A(n285), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U152 ( .A(n207), .B(B[16]), .Z(DIFF[16]) );
  NAND3_X1 U153 ( .A1(n224), .A2(n225), .A3(n289), .ZN(n287) );
  XOR2_X1 U155 ( .A(n291), .B(B[12]), .Z(DIFF[12]) );
  XOR2_X1 U156 ( .A(n294), .B(B[10]), .Z(DIFF[10]) );
  NAND3_X1 U157 ( .A1(n243), .A2(n221), .A3(n295), .ZN(n234) );
  NOR3_X1 U3 ( .A1(B[30]), .A2(B[31]), .A3(n272), .ZN(n270) );
  OR2_X1 U4 ( .A1(B[26]), .A2(B[27]), .ZN(n204) );
  OR2_X1 U5 ( .A1(B[22]), .A2(B[23]), .ZN(n205) );
  OR2_X1 U6 ( .A1(B[17]), .A2(B[16]), .ZN(n206) );
  NAND3_X1 U7 ( .A1(n224), .A2(n225), .A3(n289), .ZN(n207) );
  CLKBUF_X1 U8 ( .A(n234), .Z(n208) );
  NOR2_X1 U9 ( .A1(n294), .A2(B[10]), .ZN(n209) );
  AND2_X1 U10 ( .A1(n209), .A2(n210), .ZN(n289) );
  AND2_X1 U11 ( .A1(n219), .A2(n223), .ZN(n210) );
  BUF_X1 U12 ( .A(n283), .Z(n216) );
  BUF_X1 U13 ( .A(n289), .Z(n214) );
  OR2_X1 U14 ( .A1(n234), .A2(n211), .ZN(n294) );
  OR2_X1 U15 ( .A1(B[8]), .A2(B[9]), .ZN(n211) );
  XOR2_X1 U16 ( .A(n212), .B(n225), .Z(DIFF[15]) );
  AND2_X1 U17 ( .A1(n214), .A2(n224), .ZN(n212) );
  AND2_X1 U18 ( .A1(n275), .A2(n213), .ZN(n243) );
  NOR2_X1 U19 ( .A1(B[2]), .A2(B[3]), .ZN(n213) );
  CLKBUF_X1 U20 ( .A(n279), .Z(n215) );
  NOR2_X1 U21 ( .A1(n277), .A2(n204), .ZN(n217) );
  NOR2_X1 U22 ( .A1(n277), .A2(n204), .ZN(n274) );
  NOR2_X1 U23 ( .A1(n264), .A2(B[3]), .ZN(n218) );
  NOR2_X1 U24 ( .A1(n287), .A2(n206), .ZN(n286) );
  NOR2_X1 U25 ( .A1(n281), .A2(n205), .ZN(n279) );
  NOR2_X1 U26 ( .A1(B[13]), .A2(B[12]), .ZN(n219) );
  XOR2_X1 U27 ( .A(n301), .B(n259), .Z(DIFF[43]) );
  XOR2_X1 U28 ( .A(n298), .B(n265), .Z(DIFF[38]) );
  NOR3_X1 U29 ( .A1(B[48]), .A2(B[49]), .A3(n253), .ZN(n251) );
  NOR3_X1 U30 ( .A1(B[52]), .A2(B[53]), .A3(n249), .ZN(n247) );
  NOR3_X1 U31 ( .A1(B[56]), .A2(B[57]), .A3(n245), .ZN(n242) );
  NOR3_X1 U32 ( .A1(B[44]), .A2(B[45]), .A3(n257), .ZN(n255) );
  NOR3_X1 U33 ( .A1(B[60]), .A2(B[61]), .A3(n240), .ZN(n239) );
  NOR2_X1 U34 ( .A1(n263), .A2(B[39]), .ZN(n261) );
  XOR2_X1 U35 ( .A(n297), .B(n268), .Z(DIFF[35]) );
  NOR2_X1 U36 ( .A1(n260), .A2(B[42]), .ZN(n259) );
  XNOR2_X1 U37 ( .A(B[37]), .B(n267), .ZN(DIFF[37]) );
  NOR2_X1 U38 ( .A1(n237), .A2(B[5]), .ZN(n236) );
  NOR2_X1 U39 ( .A1(n269), .A2(B[34]), .ZN(n268) );
  XNOR2_X1 U40 ( .A(n236), .B(B[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U41 ( .A(n284), .B(n228), .ZN(DIFF[21]) );
  XNOR2_X1 U42 ( .A(n280), .B(n230), .ZN(DIFF[25]) );
  NAND2_X1 U43 ( .A1(n236), .A2(n222), .ZN(n235) );
  XOR2_X1 U44 ( .A(n223), .B(n293), .Z(DIFF[11]) );
  NOR2_X1 U45 ( .A1(n285), .A2(B[19]), .ZN(n283) );
  XNOR2_X1 U46 ( .A(n276), .B(n232), .ZN(DIFF[29]) );
  NOR2_X1 U47 ( .A1(n294), .A2(B[10]), .ZN(n293) );
  XOR2_X1 U48 ( .A(n275), .B(n220), .Z(DIFF[2]) );
  XOR2_X1 U49 ( .A(n226), .B(n286), .Z(DIFF[18]) );
  XNOR2_X1 U50 ( .A(B[53]), .B(n250), .ZN(DIFF[53]) );
  NOR2_X1 U51 ( .A1(B[52]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U52 ( .A(B[50]), .B(n251), .ZN(DIFF[50]) );
  XNOR2_X1 U53 ( .A(B[45]), .B(n258), .ZN(DIFF[45]) );
  NOR2_X1 U54 ( .A1(B[44]), .A2(n257), .ZN(n258) );
  XNOR2_X1 U55 ( .A(B[46]), .B(n255), .ZN(DIFF[46]) );
  XNOR2_X1 U56 ( .A(B[54]), .B(n247), .ZN(DIFF[54]) );
  NAND2_X1 U57 ( .A1(n251), .A2(n304), .ZN(n252) );
  NAND2_X1 U58 ( .A1(n255), .A2(n302), .ZN(n256) );
  NAND2_X1 U59 ( .A1(n247), .A2(n306), .ZN(n248) );
  XNOR2_X1 U60 ( .A(B[57]), .B(n246), .ZN(DIFF[57]) );
  NOR2_X1 U61 ( .A1(B[56]), .A2(n245), .ZN(n246) );
  NAND2_X1 U62 ( .A1(n239), .A2(n310), .ZN(n238) );
  XNOR2_X1 U63 ( .A(B[61]), .B(n241), .ZN(DIFF[61]) );
  NOR2_X1 U64 ( .A1(B[60]), .A2(n240), .ZN(n241) );
  XNOR2_X1 U65 ( .A(B[62]), .B(n239), .ZN(DIFF[62]) );
  NAND2_X1 U66 ( .A1(n242), .A2(n308), .ZN(n244) );
  XNOR2_X1 U67 ( .A(B[58]), .B(n242), .ZN(DIFF[58]) );
  XNOR2_X1 U68 ( .A(n271), .B(n296), .ZN(DIFF[33]) );
  XNOR2_X1 U69 ( .A(B[13]), .B(n292), .ZN(DIFF[13]) );
  XNOR2_X1 U70 ( .A(B[32]), .B(n270), .ZN(DIFF[32]) );
  XNOR2_X1 U71 ( .A(B[49]), .B(n254), .ZN(DIFF[49]) );
  NOR2_X1 U72 ( .A1(B[48]), .A2(n253), .ZN(n254) );
  NOR2_X1 U73 ( .A1(B[1]), .A2(\B[0] ), .ZN(n275) );
  NOR3_X1 U74 ( .A1(B[7]), .A2(B[5]), .A3(B[6]), .ZN(n295) );
  NAND2_X1 U75 ( .A1(n218), .A2(n221), .ZN(n237) );
  XNOR2_X1 U76 ( .A(n243), .B(B[4]), .ZN(DIFF[4]) );
  NAND2_X1 U77 ( .A1(n215), .A2(n229), .ZN(n280) );
  XNOR2_X1 U78 ( .A(B[24]), .B(n215), .ZN(DIFF[24]) );
  XNOR2_X1 U79 ( .A(B[17]), .B(n288), .ZN(DIFF[17]) );
  NAND2_X1 U80 ( .A1(n259), .A2(n301), .ZN(n257) );
  NAND2_X1 U81 ( .A1(n261), .A2(n299), .ZN(n262) );
  XNOR2_X1 U82 ( .A(B[40]), .B(n261), .ZN(DIFF[40]) );
  XNOR2_X1 U83 ( .A(B[31]), .B(n273), .ZN(DIFF[31]) );
  OR2_X1 U84 ( .A1(n234), .A2(B[8]), .ZN(n233) );
  NAND2_X1 U85 ( .A1(n270), .A2(n290), .ZN(n271) );
  XNOR2_X1 U86 ( .A(B[27]), .B(n278), .ZN(DIFF[27]) );
  NOR2_X1 U87 ( .A1(B[12]), .A2(n291), .ZN(n292) );
  NOR2_X1 U88 ( .A1(B[36]), .A2(n266), .ZN(n267) );
  NOR3_X1 U89 ( .A1(B[36]), .A2(B[37]), .A3(n266), .ZN(n265) );
  XNOR2_X1 U90 ( .A(B[23]), .B(n282), .ZN(DIFF[23]) );
  NAND2_X1 U91 ( .A1(n293), .A2(n223), .ZN(n291) );
  NAND2_X1 U92 ( .A1(n265), .A2(n298), .ZN(n263) );
  NAND2_X1 U93 ( .A1(n275), .A2(n220), .ZN(n264) );
  XNOR2_X1 U94 ( .A(B[20]), .B(n216), .ZN(DIFF[20]) );
  NOR2_X1 U95 ( .A1(B[22]), .A2(n281), .ZN(n282) );
  NAND2_X1 U96 ( .A1(n216), .A2(n227), .ZN(n284) );
  NOR2_X1 U97 ( .A1(B[26]), .A2(n277), .ZN(n278) );
  XNOR2_X1 U98 ( .A(B[28]), .B(n217), .ZN(DIFF[28]) );
  NOR2_X1 U99 ( .A1(B[30]), .A2(n272), .ZN(n273) );
  NAND2_X1 U100 ( .A1(n217), .A2(n231), .ZN(n276) );
  NOR2_X1 U101 ( .A1(B[16]), .A2(n207), .ZN(n288) );
  XNOR2_X1 U102 ( .A(n214), .B(B[14]), .ZN(DIFF[14]) );
  NAND2_X1 U103 ( .A1(n268), .A2(n297), .ZN(n266) );
  NAND2_X1 U104 ( .A1(n286), .A2(n226), .ZN(n285) );
  INV_X1 U105 ( .A(B[2]), .ZN(n220) );
  INV_X1 U106 ( .A(B[4]), .ZN(n221) );
  INV_X1 U107 ( .A(B[6]), .ZN(n222) );
  INV_X1 U108 ( .A(B[11]), .ZN(n223) );
  INV_X1 U109 ( .A(B[14]), .ZN(n224) );
  INV_X1 U110 ( .A(B[15]), .ZN(n225) );
  INV_X1 U111 ( .A(B[18]), .ZN(n226) );
  INV_X1 U112 ( .A(B[20]), .ZN(n227) );
  INV_X1 U113 ( .A(B[21]), .ZN(n228) );
  INV_X1 U140 ( .A(B[24]), .ZN(n229) );
  INV_X1 U143 ( .A(B[25]), .ZN(n230) );
  INV_X1 U146 ( .A(B[28]), .ZN(n231) );
  INV_X1 U149 ( .A(B[29]), .ZN(n232) );
  INV_X1 U154 ( .A(B[32]), .ZN(n290) );
  INV_X1 U158 ( .A(B[33]), .ZN(n296) );
  INV_X1 U159 ( .A(B[35]), .ZN(n297) );
  INV_X1 U160 ( .A(B[38]), .ZN(n298) );
  INV_X1 U161 ( .A(B[40]), .ZN(n299) );
  INV_X1 U162 ( .A(B[41]), .ZN(n300) );
  INV_X1 U163 ( .A(B[43]), .ZN(n301) );
  INV_X1 U164 ( .A(B[46]), .ZN(n302) );
  INV_X1 U165 ( .A(B[47]), .ZN(n303) );
  INV_X1 U166 ( .A(B[50]), .ZN(n304) );
  INV_X1 U167 ( .A(B[51]), .ZN(n305) );
  INV_X1 U168 ( .A(B[54]), .ZN(n306) );
  INV_X1 U169 ( .A(B[55]), .ZN(n307) );
  INV_X1 U170 ( .A(B[58]), .ZN(n308) );
  INV_X1 U171 ( .A(B[59]), .ZN(n309) );
  INV_X1 U172 ( .A(B[62]), .ZN(n310) );
endmodule


module complement_NBIT64_30 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_30_DW01_sub_4 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_29_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n239, n240, n241, n243, n244, n245, n247, n248, n249, n251,
         n252, n253, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n238, n242, n246, n250, n254, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U114 ( .A(B[9]), .B(n227), .Z(DIFF[9]) );
  XOR2_X1 U115 ( .A(n228), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U116 ( .A(n229), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U117 ( .A(n232), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U118 ( .A(n234), .B(B[60]), .Z(DIFF[60]) );
  NAND3_X1 U119 ( .A1(n304), .A2(n305), .A3(n236), .ZN(n234) );
  XOR2_X1 U120 ( .A(n231), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U122 ( .A(n239), .B(B[56]), .Z(DIFF[56]) );
  NAND3_X1 U123 ( .A1(n302), .A2(n303), .A3(n241), .ZN(n239) );
  XOR2_X1 U125 ( .A(n243), .B(B[52]), .Z(DIFF[52]) );
  NAND3_X1 U126 ( .A1(n300), .A2(n301), .A3(n245), .ZN(n243) );
  XOR2_X1 U128 ( .A(n247), .B(B[48]), .Z(DIFF[48]) );
  NAND3_X1 U129 ( .A1(n298), .A2(n299), .A3(n249), .ZN(n247) );
  XOR2_X1 U131 ( .A(n251), .B(B[44]), .Z(DIFF[44]) );
  NAND3_X1 U132 ( .A1(n296), .A2(n297), .A3(n253), .ZN(n251) );
  XOR2_X1 U134 ( .A(n255), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U135 ( .A(n258), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U136 ( .A(n259), .B(B[38]), .Z(DIFF[38]) );
  NAND3_X1 U137 ( .A1(n292), .A2(n294), .A3(n260), .ZN(n259) );
  XOR2_X1 U138 ( .A(n261), .B(n293), .Z(DIFF[37]) );
  XOR2_X1 U139 ( .A(n262), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U140 ( .A(n264), .B(B[32]), .Z(DIFF[32]) );
  NAND3_X1 U141 ( .A1(n250), .A2(n254), .A3(n266), .ZN(n264) );
  XOR2_X1 U143 ( .A(n268), .B(B[28]), .Z(DIFF[28]) );
  XOR2_X1 U146 ( .A(n273), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U149 ( .A(n277), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U150 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U151 ( .A(n280), .B(B[18]), .Z(DIFF[18]) );
  NAND3_X1 U152 ( .A1(n223), .A2(n224), .A3(n281), .ZN(n280) );
  XOR2_X1 U154 ( .A(n205), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U155 ( .A(n286), .B(B[12]), .Z(DIFF[12]) );
  XOR2_X1 U156 ( .A(n288), .B(B[10]), .Z(DIFF[10]) );
  NAND3_X1 U157 ( .A1(n289), .A2(n218), .A3(n237), .ZN(n228) );
  NOR2_X1 U3 ( .A1(n273), .A2(n199), .ZN(n271) );
  NOR3_X1 U4 ( .A1(B[40]), .A2(B[41]), .A3(n255), .ZN(n253) );
  NOR3_X1 U5 ( .A1(B[44]), .A2(B[45]), .A3(n251), .ZN(n249) );
  OR2_X1 U6 ( .A1(B[14]), .A2(B[15]), .ZN(n198) );
  OR2_X1 U7 ( .A1(B[24]), .A2(B[25]), .ZN(n199) );
  OR2_X1 U8 ( .A1(B[20]), .A2(B[21]), .ZN(n200) );
  OR2_X1 U9 ( .A1(B[28]), .A2(B[29]), .ZN(n201) );
  AND2_X1 U10 ( .A1(n226), .A2(n238), .ZN(n202) );
  AND2_X1 U11 ( .A1(n242), .A2(n246), .ZN(n203) );
  NAND2_X1 U12 ( .A1(n210), .A2(n221), .ZN(n204) );
  NAND2_X1 U13 ( .A1(n285), .A2(n222), .ZN(n205) );
  OR2_X2 U14 ( .A1(n228), .A2(n206), .ZN(n288) );
  OR2_X1 U15 ( .A1(B[8]), .A2(B[9]), .ZN(n206) );
  NOR2_X2 U16 ( .A1(n288), .A2(n207), .ZN(n285) );
  OR2_X1 U17 ( .A1(B[10]), .A2(n204), .ZN(n207) );
  NOR2_X1 U18 ( .A1(n277), .A2(n200), .ZN(n208) );
  OR2_X1 U19 ( .A1(n280), .A2(n209), .ZN(n277) );
  OR2_X1 U20 ( .A1(B[18]), .A2(B[19]), .ZN(n209) );
  INV_X1 U21 ( .A(B[12]), .ZN(n210) );
  NOR2_X1 U22 ( .A1(n283), .A2(n198), .ZN(n211) );
  NAND2_X1 U23 ( .A1(n275), .A2(n202), .ZN(n273) );
  NAND2_X1 U24 ( .A1(n271), .A2(n203), .ZN(n268) );
  NOR2_X1 U25 ( .A1(n268), .A2(n201), .ZN(n266) );
  XNOR2_X1 U26 ( .A(n212), .B(n299), .ZN(DIFF[47]) );
  NAND2_X1 U27 ( .A1(n249), .A2(n298), .ZN(n212) );
  XNOR2_X1 U28 ( .A(n213), .B(n303), .ZN(DIFF[55]) );
  NAND2_X1 U29 ( .A1(n241), .A2(n302), .ZN(n213) );
  XNOR2_X1 U30 ( .A(n214), .B(n301), .ZN(DIFF[51]) );
  NAND2_X1 U31 ( .A1(n245), .A2(n300), .ZN(n214) );
  XNOR2_X1 U32 ( .A(n215), .B(n305), .ZN(DIFF[59]) );
  NAND2_X1 U33 ( .A1(n236), .A2(n304), .ZN(n215) );
  XOR2_X1 U34 ( .A(n216), .B(n297), .Z(DIFF[43]) );
  AND2_X1 U35 ( .A1(n253), .A2(n296), .ZN(n216) );
  OR2_X1 U36 ( .A1(B[33]), .A2(B[32]), .ZN(n217) );
  NOR2_X1 U37 ( .A1(n283), .A2(n198), .ZN(n281) );
  NOR2_X1 U38 ( .A1(n277), .A2(n200), .ZN(n275) );
  NOR2_X1 U39 ( .A1(n264), .A2(n217), .ZN(n263) );
  XOR2_X1 U40 ( .A(n295), .B(n257), .Z(DIFF[39]) );
  XOR2_X1 U41 ( .A(n306), .B(n233), .Z(DIFF[62]) );
  NOR3_X1 U42 ( .A1(B[48]), .A2(B[49]), .A3(n247), .ZN(n245) );
  NOR3_X1 U43 ( .A1(B[52]), .A2(B[53]), .A3(n243), .ZN(n241) );
  NOR3_X1 U44 ( .A1(B[56]), .A2(B[57]), .A3(n239), .ZN(n236) );
  NOR3_X1 U45 ( .A1(B[60]), .A2(B[61]), .A3(n234), .ZN(n233) );
  NAND2_X1 U46 ( .A1(n233), .A2(n306), .ZN(n232) );
  NOR2_X1 U47 ( .A1(n259), .A2(B[38]), .ZN(n257) );
  XNOR2_X1 U48 ( .A(B[41]), .B(n256), .ZN(DIFF[41]) );
  NOR2_X1 U49 ( .A1(B[40]), .A2(n255), .ZN(n256) );
  XNOR2_X1 U50 ( .A(B[49]), .B(n248), .ZN(DIFF[49]) );
  NOR2_X1 U51 ( .A1(B[48]), .A2(n247), .ZN(n248) );
  XNOR2_X1 U52 ( .A(B[53]), .B(n244), .ZN(DIFF[53]) );
  NOR2_X1 U53 ( .A1(B[52]), .A2(n243), .ZN(n244) );
  XNOR2_X1 U54 ( .A(B[45]), .B(n252), .ZN(DIFF[45]) );
  NOR2_X1 U55 ( .A1(B[44]), .A2(n251), .ZN(n252) );
  XNOR2_X1 U56 ( .A(B[57]), .B(n240), .ZN(DIFF[57]) );
  NOR2_X1 U57 ( .A1(B[56]), .A2(n239), .ZN(n240) );
  XNOR2_X1 U58 ( .A(B[61]), .B(n235), .ZN(DIFF[61]) );
  NOR2_X1 U59 ( .A1(B[60]), .A2(n234), .ZN(n235) );
  XNOR2_X1 U60 ( .A(B[50]), .B(n245), .ZN(DIFF[50]) );
  XNOR2_X1 U61 ( .A(B[54]), .B(n241), .ZN(DIFF[54]) );
  XNOR2_X1 U62 ( .A(B[46]), .B(n249), .ZN(DIFF[46]) );
  XNOR2_X1 U63 ( .A(B[58]), .B(n236), .ZN(DIFF[58]) );
  NOR2_X1 U64 ( .A1(n262), .A2(B[35]), .ZN(n260) );
  NOR2_X1 U65 ( .A1(n231), .A2(B[5]), .ZN(n230) );
  XNOR2_X1 U66 ( .A(n230), .B(n219), .ZN(DIFF[6]) );
  XNOR2_X1 U67 ( .A(n276), .B(n238), .ZN(DIFF[23]) );
  XNOR2_X1 U68 ( .A(n272), .B(n246), .ZN(DIFF[27]) );
  XOR2_X1 U69 ( .A(n222), .B(n285), .Z(DIFF[13]) );
  XOR2_X1 U70 ( .A(n225), .B(n279), .Z(DIFF[19]) );
  NAND2_X1 U71 ( .A1(n237), .A2(n218), .ZN(n231) );
  XNOR2_X1 U72 ( .A(B[25]), .B(n274), .ZN(DIFF[25]) );
  XNOR2_X1 U73 ( .A(B[21]), .B(n278), .ZN(DIFF[21]) );
  XNOR2_X1 U74 ( .A(n282), .B(n224), .ZN(DIFF[17]) );
  XNOR2_X1 U75 ( .A(n267), .B(n254), .ZN(DIFF[31]) );
  NOR2_X1 U76 ( .A1(n258), .A2(B[3]), .ZN(n237) );
  XNOR2_X1 U77 ( .A(B[29]), .B(n270), .ZN(DIFF[29]) );
  XNOR2_X1 U78 ( .A(B[33]), .B(n265), .ZN(DIFF[33]) );
  NOR2_X1 U79 ( .A1(n288), .A2(B[10]), .ZN(n287) );
  XNOR2_X1 U80 ( .A(n269), .B(B[2]), .ZN(DIFF[2]) );
  NAND2_X1 U81 ( .A1(n269), .A2(n307), .ZN(n258) );
  INV_X1 U82 ( .A(B[2]), .ZN(n307) );
  NOR2_X1 U83 ( .A1(B[1]), .A2(\B[0] ), .ZN(n269) );
  XNOR2_X1 U84 ( .A(B[42]), .B(n253), .ZN(DIFF[42]) );
  NAND2_X1 U85 ( .A1(n230), .A2(n220), .ZN(n229) );
  NAND2_X1 U86 ( .A1(n257), .A2(n295), .ZN(n255) );
  XNOR2_X1 U87 ( .A(B[15]), .B(n284), .ZN(DIFF[15]) );
  XNOR2_X1 U88 ( .A(B[36]), .B(n260), .ZN(DIFF[36]) );
  NAND2_X1 U89 ( .A1(n260), .A2(n292), .ZN(n261) );
  NOR2_X1 U90 ( .A1(B[32]), .A2(n264), .ZN(n265) );
  NOR2_X1 U91 ( .A1(B[28]), .A2(n268), .ZN(n270) );
  NOR2_X1 U92 ( .A1(B[20]), .A2(n277), .ZN(n278) );
  NOR2_X1 U93 ( .A1(n280), .A2(B[18]), .ZN(n279) );
  NOR2_X1 U94 ( .A1(B[14]), .A2(n205), .ZN(n284) );
  XNOR2_X1 U95 ( .A(B[11]), .B(n287), .ZN(DIFF[11]) );
  NAND2_X1 U96 ( .A1(n285), .A2(n222), .ZN(n283) );
  NAND2_X1 U97 ( .A1(n287), .A2(n221), .ZN(n286) );
  XNOR2_X1 U98 ( .A(n290), .B(n263), .ZN(DIFF[34]) );
  NAND2_X1 U99 ( .A1(n263), .A2(n291), .ZN(n262) );
  NOR2_X1 U100 ( .A1(B[24]), .A2(n273), .ZN(n274) );
  XNOR2_X1 U101 ( .A(n237), .B(B[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U102 ( .A(B[30]), .B(n266), .ZN(DIFF[30]) );
  NAND2_X1 U103 ( .A1(n266), .A2(n250), .ZN(n267) );
  XNOR2_X1 U104 ( .A(B[26]), .B(n271), .ZN(DIFF[26]) );
  NAND2_X1 U105 ( .A1(n271), .A2(n242), .ZN(n272) );
  XNOR2_X1 U106 ( .A(B[22]), .B(n208), .ZN(DIFF[22]) );
  NAND2_X1 U107 ( .A1(n208), .A2(n226), .ZN(n276) );
  NAND2_X1 U108 ( .A1(n211), .A2(n223), .ZN(n282) );
  XNOR2_X1 U109 ( .A(B[16]), .B(n211), .ZN(DIFF[16]) );
  OR2_X1 U110 ( .A1(n228), .A2(B[8]), .ZN(n227) );
  NOR3_X1 U111 ( .A1(B[5]), .A2(B[7]), .A3(n219), .ZN(n289) );
  INV_X1 U112 ( .A(B[4]), .ZN(n218) );
  INV_X1 U113 ( .A(n220), .ZN(n219) );
  INV_X1 U121 ( .A(B[6]), .ZN(n220) );
  INV_X1 U124 ( .A(B[11]), .ZN(n221) );
  INV_X1 U127 ( .A(B[13]), .ZN(n222) );
  INV_X1 U130 ( .A(B[16]), .ZN(n223) );
  INV_X1 U133 ( .A(B[17]), .ZN(n224) );
  INV_X1 U142 ( .A(B[19]), .ZN(n225) );
  INV_X1 U144 ( .A(B[22]), .ZN(n226) );
  INV_X1 U145 ( .A(B[23]), .ZN(n238) );
  INV_X1 U147 ( .A(B[26]), .ZN(n242) );
  INV_X1 U148 ( .A(B[27]), .ZN(n246) );
  INV_X1 U153 ( .A(B[30]), .ZN(n250) );
  INV_X1 U158 ( .A(B[31]), .ZN(n254) );
  INV_X1 U159 ( .A(n291), .ZN(n290) );
  INV_X1 U160 ( .A(B[34]), .ZN(n291) );
  INV_X1 U161 ( .A(B[36]), .ZN(n292) );
  INV_X1 U162 ( .A(n294), .ZN(n293) );
  INV_X1 U163 ( .A(B[37]), .ZN(n294) );
  INV_X1 U164 ( .A(B[39]), .ZN(n295) );
  INV_X1 U165 ( .A(B[42]), .ZN(n296) );
  INV_X1 U166 ( .A(B[43]), .ZN(n297) );
  INV_X1 U167 ( .A(B[46]), .ZN(n298) );
  INV_X1 U168 ( .A(B[47]), .ZN(n299) );
  INV_X1 U169 ( .A(B[50]), .ZN(n300) );
  INV_X1 U170 ( .A(B[51]), .ZN(n301) );
  INV_X1 U171 ( .A(B[54]), .ZN(n302) );
  INV_X1 U172 ( .A(B[55]), .ZN(n303) );
  INV_X1 U173 ( .A(B[58]), .ZN(n304) );
  INV_X1 U174 ( .A(B[59]), .ZN(n305) );
  INV_X1 U175 ( .A(B[62]), .ZN(n306) );
endmodule


module complement_NBIT64_29 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_29_DW01_sub_4 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_28_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n214, n215, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n253, n254, n255, n256, n257, n258,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n216, n252, n259, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U97 ( .A(B[9]), .B(n214), .Z(DIFF[9]) );
  XOR2_X1 U99 ( .A(n217), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U100 ( .A(n218), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U101 ( .A(n220), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U102 ( .A(n223), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U103 ( .A(n224), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U104 ( .A(n222), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U105 ( .A(n225), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U106 ( .A(n228), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U107 ( .A(n227), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U108 ( .A(n229), .B(B[52]), .Z(DIFF[52]) );
  XOR2_X1 U109 ( .A(n232), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U110 ( .A(n231), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U111 ( .A(n233), .B(B[48]), .Z(DIFF[48]) );
  XOR2_X1 U112 ( .A(n237), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U113 ( .A(n236), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U114 ( .A(n238), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U115 ( .A(n241), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U116 ( .A(n240), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U117 ( .A(n242), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U118 ( .A(n245), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U120 ( .A(n248), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U121 ( .A(n247), .B(B[36]), .Z(DIFF[36]) );
  XOR2_X1 U122 ( .A(n249), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U123 ( .A(n251), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U124 ( .A(n254), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U125 ( .A(n253), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U126 ( .A(n255), .B(B[28]), .Z(DIFF[28]) );
  XOR2_X1 U129 ( .A(n260), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U130 ( .A(n263), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U131 ( .A(n262), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U132 ( .A(n265), .B(B[20]), .Z(DIFF[20]) );
  NAND3_X1 U133 ( .A1(n266), .A2(n280), .A3(n267), .ZN(n265) );
  XOR2_X1 U134 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U135 ( .A(n268), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U136 ( .A(n272), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U137 ( .A(n271), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U138 ( .A(n273), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U139 ( .A(n275), .B(B[10]), .Z(DIFF[10]) );
  OR2_X1 U3 ( .A1(n223), .A2(B[5]), .ZN(n217) );
  NOR2_X1 U4 ( .A1(n246), .A2(B[38]), .ZN(n244) );
  NOR3_X1 U5 ( .A1(B[6]), .A2(B[7]), .A3(n217), .ZN(n215) );
  OR2_X1 U6 ( .A1(n273), .A2(B[13]), .ZN(n271) );
  INV_X1 U7 ( .A(B[27]), .ZN(n211) );
  INV_X1 U8 ( .A(B[26]), .ZN(n208) );
  NOR3_X1 U9 ( .A1(B[32]), .A2(B[33]), .A3(n251), .ZN(n250) );
  OR2_X1 U10 ( .A1(n210), .A2(n242), .ZN(n240) );
  INV_X1 U11 ( .A(B[38]), .ZN(n209) );
  OR3_X1 U12 ( .A1(B[44]), .A2(B[45]), .A3(n238), .ZN(n236) );
  OR3_X1 U13 ( .A1(B[48]), .A2(B[49]), .A3(n233), .ZN(n231) );
  OR2_X1 U14 ( .A1(B[15]), .A2(B[14]), .ZN(n203) );
  NOR3_X1 U15 ( .A1(B[10]), .A2(B[11]), .A3(n275), .ZN(n204) );
  NOR3_X1 U16 ( .A1(B[10]), .A2(B[11]), .A3(n275), .ZN(n274) );
  NAND2_X1 U17 ( .A1(n274), .A2(n279), .ZN(n205) );
  NOR2_X1 U18 ( .A1(n205), .A2(n206), .ZN(n266) );
  OR2_X1 U19 ( .A1(n203), .A2(B[13]), .ZN(n206) );
  XOR2_X1 U20 ( .A(n207), .B(n211), .Z(DIFF[27]) );
  NOR2_X1 U21 ( .A1(n258), .A2(B[26]), .ZN(n207) );
  XNOR2_X1 U22 ( .A(n258), .B(n208), .ZN(DIFF[26]) );
  XNOR2_X1 U23 ( .A(n246), .B(n209), .ZN(DIFF[38]) );
  OR2_X1 U24 ( .A1(B[41]), .A2(B[40]), .ZN(n210) );
  OR2_X1 U25 ( .A1(B[29]), .A2(B[28]), .ZN(n212) );
  OR2_X2 U26 ( .A1(n212), .A2(n255), .ZN(n253) );
  OR2_X1 U27 ( .A1(B[26]), .A2(B[27]), .ZN(n213) );
  OR2_X2 U28 ( .A1(n213), .A2(n258), .ZN(n255) );
  OR2_X2 U29 ( .A1(n214), .A2(B[9]), .ZN(n275) );
  OR3_X2 U30 ( .A1(B[36]), .A2(B[37]), .A3(n247), .ZN(n246) );
  OR3_X2 U31 ( .A1(B[24]), .A2(B[25]), .A3(n260), .ZN(n258) );
  OR3_X2 U32 ( .A1(B[30]), .A2(B[31]), .A3(n253), .ZN(n251) );
  XOR2_X1 U33 ( .A(B[33]), .B(n216), .Z(DIFF[33]) );
  OR2_X1 U34 ( .A1(B[32]), .A2(n251), .ZN(n216) );
  NAND2_X1 U35 ( .A1(n244), .A2(n285), .ZN(n242) );
  NOR3_X1 U36 ( .A1(B[60]), .A2(B[61]), .A3(n220), .ZN(n219) );
  OR3_X1 U37 ( .A1(B[58]), .A2(B[59]), .A3(n222), .ZN(n220) );
  OR3_X1 U38 ( .A1(B[42]), .A2(B[43]), .A3(n240), .ZN(n238) );
  OR3_X1 U39 ( .A1(B[46]), .A2(B[47]), .A3(n236), .ZN(n233) );
  OR3_X1 U40 ( .A1(B[50]), .A2(B[51]), .A3(n231), .ZN(n229) );
  OR3_X1 U41 ( .A1(B[54]), .A2(B[55]), .A3(n227), .ZN(n225) );
  OR3_X1 U42 ( .A1(B[52]), .A2(B[53]), .A3(n229), .ZN(n227) );
  OR3_X1 U43 ( .A1(B[56]), .A2(B[57]), .A3(n225), .ZN(n222) );
  NAND2_X1 U44 ( .A1(n215), .A2(n278), .ZN(n214) );
  OR2_X1 U45 ( .A1(n249), .A2(B[35]), .ZN(n247) );
  XNOR2_X1 U46 ( .A(n252), .B(B[7]), .ZN(DIFF[7]) );
  NOR2_X1 U47 ( .A1(n217), .A2(B[6]), .ZN(n252) );
  NAND2_X1 U48 ( .A1(n264), .A2(n282), .ZN(n262) );
  NAND2_X1 U49 ( .A1(n204), .A2(n279), .ZN(n273) );
  NAND2_X1 U50 ( .A1(n250), .A2(n284), .ZN(n249) );
  INV_X1 U51 ( .A(n266), .ZN(n287) );
  NOR3_X1 U52 ( .A1(B[16]), .A2(B[17]), .A3(n287), .ZN(n269) );
  NOR3_X1 U53 ( .A1(B[17]), .A2(B[19]), .A3(B[18]), .ZN(n267) );
  NOR2_X1 U54 ( .A1(n265), .A2(B[20]), .ZN(n264) );
  XNOR2_X1 U55 ( .A(B[11]), .B(n276), .ZN(DIFF[11]) );
  NOR2_X1 U56 ( .A1(B[10]), .A2(n275), .ZN(n276) );
  OR3_X2 U57 ( .A1(B[22]), .A2(B[23]), .A3(n262), .ZN(n260) );
  NAND2_X1 U58 ( .A1(n234), .A2(n259), .ZN(n223) );
  OR2_X1 U59 ( .A1(n240), .A2(B[42]), .ZN(n241) );
  OR2_X1 U60 ( .A1(n236), .A2(B[46]), .ZN(n237) );
  XNOR2_X1 U61 ( .A(n250), .B(n283), .ZN(DIFF[34]) );
  XNOR2_X1 U62 ( .A(B[18]), .B(n269), .ZN(DIFF[18]) );
  NAND2_X1 U63 ( .A1(n269), .A2(n281), .ZN(n268) );
  XNOR2_X1 U64 ( .A(B[49]), .B(n235), .ZN(DIFF[49]) );
  NOR2_X1 U65 ( .A1(B[48]), .A2(n233), .ZN(n235) );
  XNOR2_X1 U66 ( .A(n264), .B(B[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U67 ( .A(B[53]), .B(n230), .ZN(DIFF[53]) );
  NOR2_X1 U68 ( .A1(B[52]), .A2(n229), .ZN(n230) );
  XNOR2_X1 U69 ( .A(B[39]), .B(n244), .ZN(DIFF[39]) );
  XNOR2_X1 U70 ( .A(B[25]), .B(n261), .ZN(DIFF[25]) );
  NOR2_X1 U71 ( .A1(B[24]), .A2(n260), .ZN(n261) );
  OR2_X1 U72 ( .A1(n231), .A2(B[50]), .ZN(n232) );
  XNOR2_X1 U73 ( .A(n234), .B(B[4]), .ZN(DIFF[4]) );
  OR2_X1 U74 ( .A1(n262), .A2(B[22]), .ZN(n263) );
  OR2_X1 U75 ( .A1(n271), .A2(B[14]), .ZN(n272) );
  XNOR2_X1 U76 ( .A(n204), .B(B[12]), .ZN(DIFF[12]) );
  OR2_X1 U77 ( .A1(n227), .A2(B[54]), .ZN(n228) );
  XNOR2_X1 U78 ( .A(B[57]), .B(n226), .ZN(DIFF[57]) );
  NOR2_X1 U79 ( .A1(B[56]), .A2(n225), .ZN(n226) );
  OR2_X1 U80 ( .A1(n222), .A2(B[58]), .ZN(n224) );
  XNOR2_X1 U81 ( .A(B[61]), .B(n221), .ZN(DIFF[61]) );
  NOR2_X1 U82 ( .A1(B[60]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U83 ( .A(n219), .B(B[62]), .ZN(DIFF[62]) );
  NAND2_X1 U84 ( .A1(n219), .A2(n286), .ZN(n218) );
  XNOR2_X1 U85 ( .A(n215), .B(n277), .ZN(DIFF[8]) );
  XNOR2_X1 U86 ( .A(B[41]), .B(n243), .ZN(DIFF[41]) );
  NOR2_X1 U87 ( .A1(B[40]), .A2(n242), .ZN(n243) );
  XNOR2_X1 U88 ( .A(B[17]), .B(n270), .ZN(DIFF[17]) );
  NOR2_X1 U89 ( .A1(B[16]), .A2(n287), .ZN(n270) );
  XNOR2_X1 U90 ( .A(B[45]), .B(n239), .ZN(DIFF[45]) );
  NOR2_X1 U91 ( .A1(B[44]), .A2(n238), .ZN(n239) );
  XNOR2_X1 U92 ( .A(B[29]), .B(n257), .ZN(DIFF[29]) );
  NOR2_X1 U93 ( .A1(B[28]), .A2(n255), .ZN(n257) );
  XNOR2_X1 U94 ( .A(n266), .B(B[16]), .ZN(DIFF[16]) );
  OR2_X1 U95 ( .A1(n247), .A2(B[36]), .ZN(n248) );
  OR2_X1 U96 ( .A1(n253), .A2(B[30]), .ZN(n254) );
  NOR2_X1 U98 ( .A1(n245), .A2(B[3]), .ZN(n234) );
  XNOR2_X1 U119 ( .A(n256), .B(B[2]), .ZN(DIFF[2]) );
  NAND2_X1 U127 ( .A1(n256), .A2(n288), .ZN(n245) );
  INV_X1 U128 ( .A(B[2]), .ZN(n288) );
  NOR2_X1 U140 ( .A1(B[1]), .A2(\B[0] ), .ZN(n256) );
  INV_X1 U141 ( .A(B[4]), .ZN(n259) );
  INV_X1 U142 ( .A(n278), .ZN(n277) );
  INV_X1 U143 ( .A(B[8]), .ZN(n278) );
  INV_X1 U144 ( .A(B[12]), .ZN(n279) );
  INV_X1 U145 ( .A(B[16]), .ZN(n280) );
  INV_X1 U146 ( .A(B[18]), .ZN(n281) );
  INV_X1 U147 ( .A(B[21]), .ZN(n282) );
  INV_X1 U148 ( .A(n284), .ZN(n283) );
  INV_X1 U149 ( .A(B[34]), .ZN(n284) );
  INV_X1 U150 ( .A(B[39]), .ZN(n285) );
  INV_X1 U151 ( .A(B[62]), .ZN(n286) );
endmodule


module complement_NBIT64_28 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_28_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_27_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n263, n264, n265, n267, n268, n269, n271, n272, n273, n274, n276,
         n277, n278, n280, n281, n282, n283, n284, n285, n287, n288, n289,
         n290, n291, n293, n294, n295, n296, n298, n299, n300, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n262, n266, n270, n275, n279, n286, n292, n297, n301,
         n318;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U122 ( .A(n255), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U123 ( .A(n256), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U124 ( .A(n258), .B(B[60]), .Z(DIFF[60]) );
  NAND3_X1 U125 ( .A1(n286), .A2(n292), .A3(n260), .ZN(n258) );
  XOR2_X1 U127 ( .A(n263), .B(B[56]), .Z(DIFF[56]) );
  NAND3_X1 U128 ( .A1(n275), .A2(n279), .A3(n265), .ZN(n263) );
  XOR2_X1 U130 ( .A(n267), .B(B[52]), .Z(DIFF[52]) );
  NAND3_X1 U131 ( .A1(n266), .A2(n270), .A3(n269), .ZN(n267) );
  XOR2_X1 U133 ( .A(n272), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U134 ( .A(n271), .B(B[48]), .Z(DIFF[48]) );
  NAND3_X1 U135 ( .A1(n251), .A2(n262), .A3(n274), .ZN(n271) );
  XOR2_X1 U137 ( .A(n276), .B(B[44]), .Z(DIFF[44]) );
  NAND3_X1 U138 ( .A1(n249), .A2(n250), .A3(n278), .ZN(n276) );
  XOR2_X1 U140 ( .A(n280), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U141 ( .A(n283), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U142 ( .A(n284), .B(B[38]), .Z(DIFF[38]) );
  NAND3_X1 U143 ( .A1(n246), .A2(n247), .A3(n285), .ZN(n284) );
  XOR2_X1 U145 ( .A(n287), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U146 ( .A(n289), .B(B[32]), .Z(DIFF[32]) );
  NAND3_X1 U147 ( .A1(n243), .A2(n244), .A3(n291), .ZN(n289) );
  XOR2_X1 U149 ( .A(n293), .B(B[28]), .Z(DIFF[28]) );
  NAND3_X1 U150 ( .A1(n241), .A2(n242), .A3(n296), .ZN(n293) );
  XOR2_X1 U152 ( .A(n298), .B(B[24]), .Z(DIFF[24]) );
  NAND3_X1 U153 ( .A1(n239), .A2(n240), .A3(n300), .ZN(n298) );
  XOR2_X1 U155 ( .A(n302), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U156 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U157 ( .A(n306), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U158 ( .A(n304), .B(B[16]), .Z(DIFF[16]) );
  XOR2_X1 U159 ( .A(n311), .B(B[15]), .Z(DIFF[15]) );
  NAND3_X1 U160 ( .A1(n235), .A2(n236), .A3(n312), .ZN(n311) );
  NAND3_X1 U161 ( .A1(n254), .A2(n230), .A3(n309), .ZN(n314) );
  XOR2_X1 U162 ( .A(n315), .B(B[11]), .Z(DIFF[11]) );
  NAND3_X1 U163 ( .A1(n233), .A2(n232), .A3(n252), .ZN(n315) );
  NOR3_X1 U3 ( .A1(n272), .A2(B[4]), .A3(n317), .ZN(n253) );
  NOR3_X1 U4 ( .A1(n304), .A2(B[16]), .A3(n305), .ZN(n303) );
  NOR2_X1 U5 ( .A1(n302), .A2(B[21]), .ZN(n300) );
  NOR3_X1 U6 ( .A1(B[24]), .A2(B[25]), .A3(n298), .ZN(n296) );
  NOR2_X1 U7 ( .A1(n284), .A2(B[38]), .ZN(n282) );
  NOR2_X1 U8 ( .A1(n287), .A2(B[35]), .ZN(n285) );
  NOR3_X1 U9 ( .A1(B[32]), .A2(B[33]), .A3(n289), .ZN(n288) );
  NOR3_X1 U10 ( .A1(B[28]), .A2(B[29]), .A3(n293), .ZN(n291) );
  NOR3_X1 U11 ( .A1(B[44]), .A2(B[45]), .A3(n276), .ZN(n274) );
  XNOR2_X1 U12 ( .A(n220), .B(n250), .ZN(DIFF[43]) );
  NAND2_X1 U13 ( .A1(n278), .A2(n249), .ZN(n220) );
  XNOR2_X1 U14 ( .A(n221), .B(n270), .ZN(DIFF[51]) );
  NAND2_X1 U15 ( .A1(n269), .A2(n266), .ZN(n221) );
  XNOR2_X1 U16 ( .A(n222), .B(n262), .ZN(DIFF[47]) );
  NAND2_X1 U17 ( .A1(n274), .A2(n251), .ZN(n222) );
  XNOR2_X1 U18 ( .A(n223), .B(n279), .ZN(DIFF[55]) );
  NAND2_X1 U19 ( .A1(n265), .A2(n275), .ZN(n223) );
  XNOR2_X1 U20 ( .A(n224), .B(n292), .ZN(DIFF[59]) );
  NAND2_X1 U21 ( .A1(n260), .A2(n286), .ZN(n224) );
  XNOR2_X1 U22 ( .A(n225), .B(n242), .ZN(DIFF[27]) );
  NAND2_X1 U23 ( .A1(n296), .A2(n241), .ZN(n225) );
  XNOR2_X1 U24 ( .A(n226), .B(n247), .ZN(DIFF[37]) );
  NAND2_X1 U25 ( .A1(n285), .A2(n246), .ZN(n226) );
  XNOR2_X1 U26 ( .A(n227), .B(n244), .ZN(DIFF[31]) );
  NAND2_X1 U27 ( .A1(n291), .A2(n243), .ZN(n227) );
  XNOR2_X1 U28 ( .A(n228), .B(n240), .ZN(DIFF[23]) );
  NAND2_X1 U29 ( .A1(n300), .A2(n239), .ZN(n228) );
  OR3_X1 U30 ( .A1(B[17]), .A2(B[19]), .A3(B[18]), .ZN(n305) );
  XOR2_X1 U31 ( .A(n297), .B(n257), .Z(DIFF[62]) );
  NOR3_X1 U32 ( .A1(B[40]), .A2(B[41]), .A3(n280), .ZN(n278) );
  NOR3_X1 U33 ( .A1(B[48]), .A2(B[49]), .A3(n271), .ZN(n269) );
  NOR3_X1 U34 ( .A1(B[52]), .A2(B[53]), .A3(n267), .ZN(n265) );
  NOR3_X1 U35 ( .A1(B[56]), .A2(B[57]), .A3(n263), .ZN(n260) );
  NOR3_X1 U36 ( .A1(B[60]), .A2(B[61]), .A3(n258), .ZN(n257) );
  NAND2_X1 U37 ( .A1(n257), .A2(n297), .ZN(n256) );
  XNOR2_X1 U38 ( .A(B[45]), .B(n277), .ZN(DIFF[45]) );
  NOR2_X1 U39 ( .A1(B[44]), .A2(n276), .ZN(n277) );
  XNOR2_X1 U40 ( .A(B[41]), .B(n281), .ZN(DIFF[41]) );
  NOR2_X1 U41 ( .A1(B[40]), .A2(n280), .ZN(n281) );
  XNOR2_X1 U42 ( .A(B[57]), .B(n264), .ZN(DIFF[57]) );
  NOR2_X1 U43 ( .A1(B[56]), .A2(n263), .ZN(n264) );
  XNOR2_X1 U44 ( .A(B[61]), .B(n259), .ZN(DIFF[61]) );
  NOR2_X1 U45 ( .A1(B[60]), .A2(n258), .ZN(n259) );
  XNOR2_X1 U46 ( .A(B[42]), .B(n278), .ZN(DIFF[42]) );
  XNOR2_X1 U47 ( .A(B[46]), .B(n274), .ZN(DIFF[46]) );
  XNOR2_X1 U48 ( .A(B[50]), .B(n269), .ZN(DIFF[50]) );
  XNOR2_X1 U49 ( .A(B[54]), .B(n265), .ZN(DIFF[54]) );
  XNOR2_X1 U50 ( .A(B[49]), .B(n273), .ZN(DIFF[49]) );
  NOR2_X1 U51 ( .A1(B[48]), .A2(n271), .ZN(n273) );
  XNOR2_X1 U52 ( .A(B[53]), .B(n268), .ZN(DIFF[53]) );
  NOR2_X1 U53 ( .A1(B[52]), .A2(n267), .ZN(n268) );
  XNOR2_X1 U54 ( .A(B[58]), .B(n260), .ZN(DIFF[58]) );
  XOR2_X1 U55 ( .A(n248), .B(n282), .Z(DIFF[39]) );
  NAND2_X1 U56 ( .A1(n282), .A2(n248), .ZN(n280) );
  XNOR2_X1 U57 ( .A(n254), .B(B[7]), .ZN(DIFF[7]) );
  NOR2_X1 U58 ( .A1(n255), .A2(B[6]), .ZN(n254) );
  XNOR2_X1 U59 ( .A(n314), .B(n234), .ZN(DIFF[12]) );
  XNOR2_X1 U60 ( .A(B[26]), .B(n296), .ZN(DIFF[26]) );
  XNOR2_X1 U61 ( .A(B[36]), .B(n285), .ZN(DIFF[36]) );
  XNOR2_X1 U62 ( .A(B[22]), .B(n300), .ZN(DIFF[22]) );
  XNOR2_X1 U63 ( .A(B[25]), .B(n299), .ZN(DIFF[25]) );
  NOR2_X1 U64 ( .A1(B[24]), .A2(n298), .ZN(n299) );
  XNOR2_X1 U65 ( .A(B[18]), .B(n307), .ZN(DIFF[18]) );
  XOR2_X1 U66 ( .A(n245), .B(n288), .Z(DIFF[34]) );
  XNOR2_X1 U67 ( .A(n313), .B(n236), .ZN(DIFF[14]) );
  NAND2_X1 U68 ( .A1(n312), .A2(n235), .ZN(n313) );
  XNOR2_X1 U69 ( .A(B[13]), .B(n312), .ZN(DIFF[13]) );
  XOR2_X1 U70 ( .A(n238), .B(n303), .Z(DIFF[20]) );
  NAND2_X1 U71 ( .A1(n288), .A2(n245), .ZN(n287) );
  NAND2_X1 U72 ( .A1(n303), .A2(n238), .ZN(n302) );
  NOR4_X1 U73 ( .A1(B[10]), .A2(B[11]), .A3(B[8]), .A4(n231), .ZN(n309) );
  NOR3_X1 U74 ( .A1(B[16]), .A2(B[17]), .A3(n304), .ZN(n307) );
  NAND4_X1 U75 ( .A1(n253), .A2(n234), .A3(n309), .A4(n310), .ZN(n304) );
  NOR3_X1 U76 ( .A1(B[13]), .A2(B[15]), .A3(B[14]), .ZN(n310) );
  NOR2_X1 U77 ( .A1(n314), .A2(B[12]), .ZN(n312) );
  NOR2_X1 U78 ( .A1(n301), .A2(B[8]), .ZN(n252) );
  INV_X1 U79 ( .A(n253), .ZN(n301) );
  NAND2_X1 U80 ( .A1(n307), .A2(n237), .ZN(n306) );
  XNOR2_X1 U81 ( .A(n253), .B(B[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U82 ( .A(B[17]), .B(n308), .ZN(DIFF[17]) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(n304), .ZN(n308) );
  XNOR2_X1 U84 ( .A(B[33]), .B(n290), .ZN(DIFF[33]) );
  NOR2_X1 U85 ( .A1(B[32]), .A2(n289), .ZN(n290) );
  XNOR2_X1 U86 ( .A(B[29]), .B(n295), .ZN(DIFF[29]) );
  NOR2_X1 U87 ( .A1(B[28]), .A2(n293), .ZN(n295) );
  XNOR2_X1 U88 ( .A(B[30]), .B(n291), .ZN(DIFF[30]) );
  NAND2_X1 U89 ( .A1(n261), .A2(n229), .ZN(n255) );
  XNOR2_X1 U90 ( .A(n261), .B(B[5]), .ZN(DIFF[5]) );
  OR3_X1 U91 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n317) );
  XNOR2_X1 U92 ( .A(n316), .B(n233), .ZN(DIFF[10]) );
  NAND2_X1 U93 ( .A1(n252), .A2(n232), .ZN(n316) );
  XNOR2_X1 U94 ( .A(n231), .B(n252), .ZN(DIFF[9]) );
  NOR2_X1 U95 ( .A1(n272), .A2(B[4]), .ZN(n261) );
  XNOR2_X1 U96 ( .A(n294), .B(B[2]), .ZN(DIFF[2]) );
  OR2_X1 U97 ( .A1(n283), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U98 ( .A1(n294), .A2(n318), .ZN(n283) );
  INV_X1 U99 ( .A(B[2]), .ZN(n318) );
  NOR2_X1 U100 ( .A1(B[1]), .A2(\B[0] ), .ZN(n294) );
  INV_X1 U101 ( .A(B[5]), .ZN(n229) );
  INV_X1 U102 ( .A(B[7]), .ZN(n230) );
  INV_X1 U103 ( .A(n232), .ZN(n231) );
  INV_X1 U104 ( .A(B[9]), .ZN(n232) );
  INV_X1 U105 ( .A(B[10]), .ZN(n233) );
  INV_X1 U106 ( .A(B[12]), .ZN(n234) );
  INV_X1 U107 ( .A(B[13]), .ZN(n235) );
  INV_X1 U108 ( .A(B[14]), .ZN(n236) );
  INV_X1 U109 ( .A(B[18]), .ZN(n237) );
  INV_X1 U110 ( .A(B[20]), .ZN(n238) );
  INV_X1 U111 ( .A(B[22]), .ZN(n239) );
  INV_X1 U112 ( .A(B[23]), .ZN(n240) );
  INV_X1 U113 ( .A(B[26]), .ZN(n241) );
  INV_X1 U114 ( .A(B[27]), .ZN(n242) );
  INV_X1 U115 ( .A(B[30]), .ZN(n243) );
  INV_X1 U116 ( .A(B[31]), .ZN(n244) );
  INV_X1 U117 ( .A(B[34]), .ZN(n245) );
  INV_X1 U118 ( .A(B[36]), .ZN(n246) );
  INV_X1 U119 ( .A(B[37]), .ZN(n247) );
  INV_X1 U120 ( .A(B[39]), .ZN(n248) );
  INV_X1 U121 ( .A(B[42]), .ZN(n249) );
  INV_X1 U126 ( .A(B[43]), .ZN(n250) );
  INV_X1 U129 ( .A(B[46]), .ZN(n251) );
  INV_X1 U132 ( .A(B[47]), .ZN(n262) );
  INV_X1 U136 ( .A(B[50]), .ZN(n266) );
  INV_X1 U139 ( .A(B[51]), .ZN(n270) );
  INV_X1 U144 ( .A(B[54]), .ZN(n275) );
  INV_X1 U148 ( .A(B[55]), .ZN(n279) );
  INV_X1 U151 ( .A(B[58]), .ZN(n286) );
  INV_X1 U154 ( .A(B[59]), .ZN(n292) );
  INV_X1 U164 ( .A(B[62]), .ZN(n297) );
endmodule


module complement_NBIT64_27 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_27_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_26_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n42, n44,
         n45, n46, n48, n49, n54, n56, n58, n60, n61, n65, n67, n70, n73, n74,
         n79, n82, n85, n86, n91, n94, n97, n98, n100, n101, n102, n106, n108,
         n109, n110, n112, n114, n118, n120, n130, n131, n133, n134, n135,
         n136, n139, n140, n141, n144, n145, n147, n148, n149, n152, n154,
         n155, n158, n159, n162, n163, n170, n171, n173, n174, n175, n176,
         n179, n180, n181, n184, n185, n186, n188, n189, n190, n194, n195,
         n196, n198, n203, n204, n205, n206, n207, n208, n209, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U7 ( .A(n3), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U10 ( .A(n4), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U12 ( .A(n360), .B(n5), .Z(DIFF[3]) );
  XOR2_X1 U43 ( .A(B[40]), .B(n114), .Z(DIFF[40]) );
  XOR2_X1 U46 ( .A(B[39]), .B(n130), .Z(DIFF[39]) );
  XOR2_X1 U48 ( .A(B[47]), .B(n108), .Z(DIFF[47]) );
  XOR2_X1 U58 ( .A(n342), .B(n352), .Z(DIFF[57]) );
  XOR2_X1 U63 ( .A(n334), .B(n350), .Z(DIFF[49]) );
  XOR2_X1 U64 ( .A(n91), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U65 ( .A(n338), .B(n351), .Z(DIFF[53]) );
  XOR2_X1 U66 ( .A(n79), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U70 ( .A(n67), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U94 ( .A(n196), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U95 ( .A(n7), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U96 ( .A(n2), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U102 ( .A(n159), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U123 ( .A(n299), .B(n195), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(B[15]), .B(n194), .Z(DIFF[15]) );
  XOR2_X1 U126 ( .A(n297), .B(n198), .Z(DIFF[12]) );
  XOR2_X1 U131 ( .A(B[31]), .B(n154), .Z(DIFF[31]) );
  XOR2_X1 U160 ( .A(B[23]), .B(n170), .Z(DIFF[23]) );
  XOR2_X1 U164 ( .A(B[10]), .B(n204), .Z(DIFF[10]) );
  XOR2_X1 U166 ( .A(B[27]), .B(n162), .Z(DIFF[27]) );
  XOR2_X1 U169 ( .A(B[19]), .B(n179), .Z(DIFF[19]) );
  XOR2_X1 U172 ( .A(B[11]), .B(n203), .Z(DIFF[11]) );
  XOR2_X1 U185 ( .A(B[35]), .B(n139), .Z(DIFF[35]) );
  XOR2_X1 U189 ( .A(n359), .B(n13), .Z(DIFF[2]) );
  XOR2_X1 U192 ( .A(\B[0] ), .B(B[1]), .Z(DIFF[1]) );
  XOR2_X1 U193 ( .A(B[5]), .B(n65), .Z(DIFF[5]) );
  NAND3_X1 U248 ( .A1(n343), .A2(n344), .A3(n342), .ZN(n61) );
  NAND3_X1 U250 ( .A1(n339), .A2(n340), .A3(n338), .ZN(n74) );
  NAND3_X1 U252 ( .A1(n335), .A2(n336), .A3(n334), .ZN(n86) );
  NAND3_X1 U254 ( .A1(n355), .A2(n10), .A3(n100), .ZN(n98) );
  NAND3_X1 U260 ( .A1(n354), .A2(n12), .A3(n147), .ZN(n145) );
  NAND3_X1 U269 ( .A1(n295), .A2(n294), .A3(n8), .ZN(n203) );
  XOR2_X1 U3 ( .A(n205), .B(n336), .Z(DIFF[51]) );
  XOR2_X1 U5 ( .A(n206), .B(n340), .Z(DIFF[55]) );
  XOR2_X1 U8 ( .A(n207), .B(n344), .Z(DIFF[59]) );
  XOR2_X1 U34 ( .A(n70), .B(n341), .Z(DIFF[56]) );
  XOR2_X1 U35 ( .A(n82), .B(n337), .Z(DIFF[52]) );
  XOR2_X1 U36 ( .A(n346), .B(n56), .Z(DIFF[61]) );
  XOR2_X1 U37 ( .A(n54), .B(n347), .Z(DIFF[62]) );
  XOR2_X1 U38 ( .A(n345), .B(n58), .Z(DIFF[60]) );
  XOR2_X1 U55 ( .A(n94), .B(n333), .Z(DIFF[48]) );
  XOR2_X1 U57 ( .A(n208), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U76 ( .A(n349), .B(n321), .Z(DIFF[36]) );
  XOR2_X1 U110 ( .A(n348), .B(n305), .Z(DIFF[20]) );
  INV_X1 U4 ( .A(n73), .ZN(n351) );
  INV_X1 U6 ( .A(n60), .ZN(n352) );
  AND2_X1 U9 ( .A1(n120), .A2(n326), .ZN(n118) );
  AND2_X1 U11 ( .A1(n110), .A2(n330), .ZN(n109) );
  AND2_X1 U13 ( .A1(n112), .A2(n329), .ZN(n110) );
  NOR2_X1 U14 ( .A1(n85), .A2(n86), .ZN(n82) );
  NOR2_X1 U15 ( .A1(n73), .A2(n74), .ZN(n70) );
  NAND2_X1 U16 ( .A1(n82), .A2(n337), .ZN(n73) );
  NAND2_X1 U17 ( .A1(n70), .A2(n341), .ZN(n60) );
  NOR2_X1 U18 ( .A1(n91), .A2(B[50]), .ZN(n205) );
  NOR2_X1 U19 ( .A1(n79), .A2(B[54]), .ZN(n206) );
  NOR2_X1 U20 ( .A1(n67), .A2(B[58]), .ZN(n207) );
  NAND2_X1 U21 ( .A1(n334), .A2(n350), .ZN(n91) );
  NAND2_X1 U22 ( .A1(n338), .A2(n351), .ZN(n79) );
  NAND2_X1 U23 ( .A1(n342), .A2(n352), .ZN(n67) );
  INV_X1 U24 ( .A(n85), .ZN(n350) );
  NAND2_X1 U25 ( .A1(n329), .A2(n330), .ZN(n102) );
  NOR2_X1 U26 ( .A1(n60), .A2(n61), .ZN(n58) );
  AND2_X1 U27 ( .A1(n346), .A2(n56), .ZN(n54) );
  AND2_X1 U28 ( .A1(n345), .A2(n58), .ZN(n56) );
  NAND2_X1 U29 ( .A1(n327), .A2(n118), .ZN(n3) );
  NOR2_X1 U30 ( .A1(n7), .A2(B[25]), .ZN(n163) );
  NOR2_X1 U31 ( .A1(n114), .A2(n106), .ZN(n112) );
  NOR2_X1 U32 ( .A1(B[40]), .A2(n114), .ZN(n120) );
  XNOR2_X1 U33 ( .A(B[41]), .B(n120), .ZN(DIFF[41]) );
  XNOR2_X1 U39 ( .A(n118), .B(B[42]), .ZN(DIFF[42]) );
  XNOR2_X1 U40 ( .A(n131), .B(B[38]), .ZN(DIFF[38]) );
  NAND2_X1 U41 ( .A1(n323), .A2(n131), .ZN(n130) );
  NAND2_X1 U42 ( .A1(n331), .A2(n109), .ZN(n108) );
  NAND4_X1 U44 ( .A1(n325), .A2(n328), .A3(n327), .A4(n326), .ZN(n106) );
  XNOR2_X1 U45 ( .A(B[44]), .B(n112), .ZN(DIFF[44]) );
  XNOR2_X1 U47 ( .A(B[45]), .B(n110), .ZN(DIFF[45]) );
  XNOR2_X1 U49 ( .A(n109), .B(B[46]), .ZN(DIFF[46]) );
  NAND2_X1 U50 ( .A1(n94), .A2(n333), .ZN(n85) );
  NAND2_X1 U51 ( .A1(n331), .A2(n332), .ZN(n101) );
  NAND2_X1 U52 ( .A1(n54), .A2(n347), .ZN(n208) );
  NOR2_X1 U53 ( .A1(n159), .A2(n152), .ZN(n158) );
  NOR2_X1 U54 ( .A1(n2), .A2(B[29]), .ZN(n155) );
  NOR2_X1 U56 ( .A1(n196), .A2(B[13]), .ZN(n195) );
  NOR2_X1 U59 ( .A1(n42), .A2(n188), .ZN(n198) );
  XNOR2_X1 U60 ( .A(B[37]), .B(n11), .ZN(DIFF[37]) );
  NAND2_X1 U61 ( .A1(n10), .A2(n349), .ZN(n114) );
  NAND2_X1 U62 ( .A1(n12), .A2(n348), .ZN(n159) );
  AND2_X1 U67 ( .A1(n9), .A2(n306), .ZN(n171) );
  AND2_X1 U68 ( .A1(n11), .A2(n322), .ZN(n131) );
  AND2_X1 U69 ( .A1(n181), .A2(n302), .ZN(n180) );
  INV_X1 U71 ( .A(n144), .ZN(n348) );
  INV_X1 U72 ( .A(n97), .ZN(n349) );
  INV_X1 U73 ( .A(n188), .ZN(n353) );
  OR2_X1 U74 ( .A1(B[24]), .A2(n159), .ZN(n7) );
  NOR2_X1 U75 ( .A1(n97), .A2(n98), .ZN(n94) );
  NOR2_X1 U77 ( .A1(n101), .A2(n102), .ZN(n100) );
  INV_X1 U78 ( .A(n106), .ZN(n355) );
  NOR2_X1 U79 ( .A1(n184), .A2(n185), .ZN(n173) );
  NAND2_X1 U80 ( .A1(n186), .A2(n353), .ZN(n185) );
  NAND2_X1 U81 ( .A1(n1), .A2(n209), .ZN(n184) );
  NOR2_X1 U82 ( .A1(n189), .A2(n190), .ZN(n186) );
  NOR2_X1 U83 ( .A1(n144), .A2(n145), .ZN(n133) );
  NOR2_X1 U84 ( .A1(n148), .A2(n149), .ZN(n147) );
  INV_X1 U85 ( .A(n152), .ZN(n354) );
  NAND2_X1 U86 ( .A1(n311), .A2(n163), .ZN(n162) );
  NAND2_X1 U87 ( .A1(n307), .A2(n171), .ZN(n170) );
  NAND2_X1 U88 ( .A1(n319), .A2(n140), .ZN(n139) );
  NAND4_X1 U89 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(n188) );
  NAND4_X1 U90 ( .A1(n309), .A2(n312), .A3(n311), .A4(n310), .ZN(n152) );
  XNOR2_X1 U91 ( .A(n8), .B(B[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U92 ( .A(B[21]), .B(n9), .ZN(DIFF[21]) );
  XNOR2_X1 U93 ( .A(n155), .B(B[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U97 ( .A(n163), .B(B[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U98 ( .A(B[17]), .B(n181), .ZN(DIFF[17]) );
  NAND2_X1 U99 ( .A1(n173), .A2(n174), .ZN(n144) );
  NOR2_X1 U100 ( .A1(n175), .A2(n176), .ZN(n174) );
  NAND2_X1 U101 ( .A1(n301), .A2(n304), .ZN(n175) );
  NAND2_X1 U103 ( .A1(n302), .A2(n303), .ZN(n176) );
  NAND2_X1 U104 ( .A1(n133), .A2(n134), .ZN(n97) );
  NOR2_X1 U105 ( .A1(n135), .A2(n136), .ZN(n134) );
  NAND2_X1 U106 ( .A1(n317), .A2(n320), .ZN(n135) );
  NAND2_X1 U107 ( .A1(n318), .A2(n319), .ZN(n136) );
  NAND2_X1 U108 ( .A1(n198), .A2(n297), .ZN(n196) );
  AND3_X1 U109 ( .A1(n293), .A2(n1), .A3(n209), .ZN(n8) );
  AND2_X1 U111 ( .A1(n141), .A2(n318), .ZN(n140) );
  NAND2_X1 U112 ( .A1(n209), .A2(n1), .ZN(n42) );
  NAND2_X1 U113 ( .A1(n158), .A2(n313), .ZN(n2) );
  AND2_X1 U114 ( .A1(n301), .A2(n173), .ZN(n181) );
  AND2_X1 U115 ( .A1(n317), .A2(n133), .ZN(n141) );
  AND2_X1 U116 ( .A1(n348), .A2(n305), .ZN(n9) );
  AND2_X1 U117 ( .A1(n349), .A2(n321), .ZN(n11) );
  AND4_X1 U118 ( .A1(n305), .A2(n308), .A3(n307), .A4(n306), .ZN(n12) );
  NAND2_X1 U119 ( .A1(n297), .A2(n298), .ZN(n190) );
  NAND2_X1 U120 ( .A1(n313), .A2(n314), .ZN(n149) );
  AND4_X1 U121 ( .A1(n321), .A2(n324), .A3(n323), .A4(n322), .ZN(n10) );
  NAND2_X1 U122 ( .A1(n303), .A2(n180), .ZN(n179) );
  NAND2_X1 U125 ( .A1(n315), .A2(n155), .ZN(n154) );
  XNOR2_X1 U127 ( .A(B[16]), .B(n173), .ZN(DIFF[16]) );
  XNOR2_X1 U128 ( .A(B[28]), .B(n158), .ZN(DIFF[28]) );
  XNOR2_X1 U129 ( .A(B[32]), .B(n133), .ZN(DIFF[32]) );
  XNOR2_X1 U130 ( .A(n140), .B(B[34]), .ZN(DIFF[34]) );
  XNOR2_X1 U132 ( .A(n180), .B(B[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U133 ( .A(B[33]), .B(n141), .ZN(DIFF[33]) );
  XNOR2_X1 U134 ( .A(n171), .B(B[22]), .ZN(DIFF[22]) );
  AND4_X1 U135 ( .A1(n291), .A2(n362), .A3(n363), .A4(n292), .ZN(n209) );
  NAND2_X1 U136 ( .A1(n299), .A2(n300), .ZN(n189) );
  NAND2_X1 U137 ( .A1(n357), .A2(n291), .ZN(n49) );
  NAND2_X1 U138 ( .A1(n315), .A2(n316), .ZN(n148) );
  AND4_X1 U139 ( .A1(n358), .A2(n357), .A3(n359), .A4(n360), .ZN(n1) );
  NAND2_X1 U140 ( .A1(n362), .A2(n363), .ZN(n48) );
  AND2_X1 U141 ( .A1(n358), .A2(n357), .ZN(n13) );
  NAND4_X1 U142 ( .A1(n293), .A2(n294), .A3(n1), .A4(n209), .ZN(n204) );
  NAND2_X1 U143 ( .A1(n299), .A2(n195), .ZN(n194) );
  XNOR2_X1 U144 ( .A(n42), .B(n293), .ZN(DIFF[8]) );
  NAND2_X1 U145 ( .A1(n1), .A2(n361), .ZN(n4) );
  INV_X1 U146 ( .A(n48), .ZN(n361) );
  XNOR2_X1 U147 ( .A(n292), .B(n44), .ZN(DIFF[7]) );
  NAND2_X1 U148 ( .A1(n45), .A2(n46), .ZN(n44) );
  NOR3_X1 U149 ( .A1(B[2]), .A2(B[3]), .A3(B[1]), .ZN(n46) );
  NOR2_X1 U150 ( .A1(n48), .A2(n49), .ZN(n45) );
  NOR2_X1 U151 ( .A1(n356), .A2(B[2]), .ZN(n5) );
  INV_X1 U152 ( .A(n13), .ZN(n356) );
  NAND2_X1 U153 ( .A1(n362), .A2(n1), .ZN(n65) );
  XNOR2_X1 U154 ( .A(n1), .B(B[4]), .ZN(DIFF[4]) );
  INV_X1 U155 ( .A(B[4]), .ZN(n362) );
  INV_X1 U156 ( .A(\B[0] ), .ZN(n357) );
  INV_X1 U157 ( .A(B[5]), .ZN(n363) );
  INV_X1 U158 ( .A(B[3]), .ZN(n360) );
  INV_X1 U159 ( .A(B[2]), .ZN(n359) );
  INV_X1 U161 ( .A(B[1]), .ZN(n358) );
  INV_X1 U162 ( .A(B[6]), .ZN(n291) );
  INV_X1 U163 ( .A(B[7]), .ZN(n292) );
  INV_X1 U165 ( .A(B[8]), .ZN(n293) );
  INV_X1 U167 ( .A(B[9]), .ZN(n294) );
  INV_X1 U168 ( .A(B[10]), .ZN(n295) );
  INV_X1 U170 ( .A(B[11]), .ZN(n296) );
  INV_X1 U171 ( .A(B[12]), .ZN(n297) );
  INV_X1 U173 ( .A(B[13]), .ZN(n298) );
  INV_X1 U174 ( .A(B[14]), .ZN(n299) );
  INV_X1 U175 ( .A(B[15]), .ZN(n300) );
  INV_X1 U176 ( .A(B[16]), .ZN(n301) );
  INV_X1 U177 ( .A(B[17]), .ZN(n302) );
  INV_X1 U178 ( .A(B[18]), .ZN(n303) );
  INV_X1 U179 ( .A(B[19]), .ZN(n304) );
  INV_X1 U180 ( .A(B[20]), .ZN(n305) );
  INV_X1 U181 ( .A(B[21]), .ZN(n306) );
  INV_X1 U182 ( .A(B[22]), .ZN(n307) );
  INV_X1 U183 ( .A(B[23]), .ZN(n308) );
  INV_X1 U184 ( .A(B[24]), .ZN(n309) );
  INV_X1 U186 ( .A(B[25]), .ZN(n310) );
  INV_X1 U187 ( .A(B[26]), .ZN(n311) );
  INV_X1 U188 ( .A(B[27]), .ZN(n312) );
  INV_X1 U190 ( .A(B[28]), .ZN(n313) );
  INV_X1 U191 ( .A(B[29]), .ZN(n314) );
  INV_X1 U194 ( .A(B[30]), .ZN(n315) );
  INV_X1 U195 ( .A(B[31]), .ZN(n316) );
  INV_X1 U196 ( .A(B[32]), .ZN(n317) );
  INV_X1 U197 ( .A(B[33]), .ZN(n318) );
  INV_X1 U198 ( .A(B[34]), .ZN(n319) );
  INV_X1 U199 ( .A(B[35]), .ZN(n320) );
  INV_X1 U200 ( .A(B[36]), .ZN(n321) );
  INV_X1 U201 ( .A(B[37]), .ZN(n322) );
  INV_X1 U202 ( .A(B[38]), .ZN(n323) );
  INV_X1 U203 ( .A(B[39]), .ZN(n324) );
  INV_X1 U204 ( .A(B[40]), .ZN(n325) );
  INV_X1 U205 ( .A(B[41]), .ZN(n326) );
  INV_X1 U206 ( .A(B[42]), .ZN(n327) );
  INV_X1 U207 ( .A(B[43]), .ZN(n328) );
  INV_X1 U208 ( .A(B[44]), .ZN(n329) );
  INV_X1 U209 ( .A(B[45]), .ZN(n330) );
  INV_X1 U210 ( .A(B[46]), .ZN(n331) );
  INV_X1 U211 ( .A(B[47]), .ZN(n332) );
  INV_X1 U212 ( .A(B[48]), .ZN(n333) );
  INV_X1 U213 ( .A(B[49]), .ZN(n334) );
  INV_X1 U214 ( .A(B[50]), .ZN(n335) );
  INV_X1 U215 ( .A(B[51]), .ZN(n336) );
  INV_X1 U216 ( .A(B[52]), .ZN(n337) );
  INV_X1 U217 ( .A(B[53]), .ZN(n338) );
  INV_X1 U218 ( .A(B[54]), .ZN(n339) );
  INV_X1 U219 ( .A(B[55]), .ZN(n340) );
  INV_X1 U220 ( .A(B[56]), .ZN(n341) );
  INV_X1 U221 ( .A(B[57]), .ZN(n342) );
  INV_X1 U222 ( .A(B[58]), .ZN(n343) );
  INV_X1 U223 ( .A(B[59]), .ZN(n344) );
  INV_X1 U224 ( .A(B[60]), .ZN(n345) );
  INV_X1 U225 ( .A(B[61]), .ZN(n346) );
  INV_X1 U226 ( .A(B[62]), .ZN(n347) );
endmodule


module complement_NBIT64_26 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_26_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_25_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n211, n212, n214, n215, n216, n217, n218, n220, n221, n222, n223,
         n225, n226, n227, n229, n230, n231, n233, n234, n235, n237, n238,
         n239, n241, n242, n243, n244, n245, n246, n247, n248, n250, n251,
         n252, n253, n255, n256, n257, n259, n260, n261, n263, n264, n265,
         n266, n267, n269, n270, n271, n272, n273, n202, n213, n219, n224,
         n228, n232, n236, n240, n249, n254, n258, n262, n268, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299;
  assign DIFF[0] = B[0];

  XOR2_X1 U97 ( .A(n214), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U98 ( .A(n216), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U100 ( .A(n218), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U101 ( .A(n220), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U103 ( .A(n223), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U104 ( .A(n225), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U106 ( .A(n227), .B(B[52]), .Z(DIFF[52]) );
  XOR2_X1 U107 ( .A(n229), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U108 ( .A(n221), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U110 ( .A(n231), .B(B[48]), .Z(DIFF[48]) );
  XOR2_X1 U111 ( .A(n233), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U113 ( .A(n235), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U114 ( .A(n237), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U116 ( .A(n239), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U117 ( .A(n242), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U119 ( .A(n244), .B(B[36]), .Z(DIFF[36]) );
  XOR2_X1 U120 ( .A(n247), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U122 ( .A(n248), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U123 ( .A(n250), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U125 ( .A(n252), .B(B[28]), .Z(DIFF[28]) );
  XOR2_X1 U126 ( .A(n255), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U128 ( .A(n257), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U129 ( .A(n259), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U131 ( .A(n261), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U132 ( .A(B[1]), .B(B[0]), .Z(DIFF[1]) );
  XOR2_X1 U133 ( .A(n263), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U134 ( .A(n265), .B(B[16]), .Z(DIFF[16]) );
  XOR2_X1 U136 ( .A(n267), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U137 ( .A(n269), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U138 ( .A(n272), .B(B[11]), .Z(DIFF[11]) );
  NAND3_X1 U139 ( .A1(n286), .A2(n285), .A3(n211), .ZN(n272) );
  XOR2_X1 U20 ( .A(n217), .B(n295), .Z(DIFF[62]) );
  XOR2_X1 U60 ( .A(n243), .B(n293), .Z(DIFF[38]) );
  XOR2_X1 U61 ( .A(n292), .B(n246), .Z(DIFF[35]) );
  XOR2_X1 U62 ( .A(n264), .B(n288), .Z(DIFF[18]) );
  XOR2_X1 U63 ( .A(n287), .B(n270), .Z(DIFF[12]) );
  OR3_X1 U3 ( .A1(B[20]), .A2(B[21]), .A3(n261), .ZN(n259) );
  OR3_X1 U4 ( .A1(B[24]), .A2(B[25]), .A3(n257), .ZN(n255) );
  OR3_X1 U5 ( .A1(B[26]), .A2(B[27]), .A3(n255), .ZN(n252) );
  OR3_X1 U6 ( .A1(B[28]), .A2(B[29]), .A3(n252), .ZN(n250) );
  AND4_X1 U7 ( .A1(n289), .A2(n290), .A3(n296), .A4(n291), .ZN(n246) );
  OR3_X1 U8 ( .A1(B[30]), .A2(B[31]), .A3(n250), .ZN(n248) );
  OR3_X1 U9 ( .A1(B[40]), .A2(B[41]), .A3(n239), .ZN(n237) );
  OR3_X1 U10 ( .A1(B[44]), .A2(B[45]), .A3(n235), .ZN(n233) );
  OR3_X1 U11 ( .A1(B[50]), .A2(B[51]), .A3(n229), .ZN(n227) );
  NOR3_X1 U12 ( .A1(B[60]), .A2(B[61]), .A3(n218), .ZN(n217) );
  OR3_X1 U13 ( .A1(B[48]), .A2(B[49]), .A3(n231), .ZN(n229) );
  OR3_X1 U14 ( .A1(B[52]), .A2(B[53]), .A3(n227), .ZN(n225) );
  OR3_X1 U15 ( .A1(B[56]), .A2(B[57]), .A3(n223), .ZN(n220) );
  OR3_X1 U16 ( .A1(B[58]), .A2(B[59]), .A3(n220), .ZN(n218) );
  OR3_X1 U17 ( .A1(B[42]), .A2(B[43]), .A3(n237), .ZN(n235) );
  OR3_X1 U18 ( .A1(B[46]), .A2(B[47]), .A3(n233), .ZN(n231) );
  OR3_X1 U19 ( .A1(B[54]), .A2(B[55]), .A3(n225), .ZN(n223) );
  NAND2_X1 U21 ( .A1(n246), .A2(n292), .ZN(n244) );
  XNOR2_X1 U22 ( .A(n273), .B(n286), .ZN(DIFF[10]) );
  NAND2_X1 U23 ( .A1(n211), .A2(n285), .ZN(n273) );
  XNOR2_X1 U24 ( .A(B[9]), .B(n211), .ZN(DIFF[9]) );
  OR2_X1 U25 ( .A1(n241), .A2(B[39]), .ZN(n239) );
  NAND2_X1 U26 ( .A1(n264), .A2(n288), .ZN(n263) );
  NAND2_X1 U27 ( .A1(n270), .A2(n287), .ZN(n269) );
  NOR3_X1 U28 ( .A1(B[16]), .A2(B[17]), .A3(n265), .ZN(n264) );
  NOR2_X1 U29 ( .A1(n297), .A2(B[8]), .ZN(n211) );
  INV_X1 U30 ( .A(n212), .ZN(n297) );
  XNOR2_X1 U31 ( .A(n212), .B(B[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U32 ( .A(n249), .B(B[15]), .ZN(DIFF[15]) );
  NOR2_X1 U33 ( .A1(n267), .A2(B[14]), .ZN(n249) );
  OR2_X1 U34 ( .A1(n269), .A2(B[13]), .ZN(n267) );
  OR2_X1 U35 ( .A1(n263), .A2(B[19]), .ZN(n261) );
  OR3_X1 U36 ( .A1(B[22]), .A2(B[23]), .A3(n259), .ZN(n257) );
  AND3_X1 U37 ( .A1(n212), .A2(n286), .A3(n271), .ZN(n270) );
  NOR3_X1 U38 ( .A1(B[11]), .A2(B[9]), .A3(B[8]), .ZN(n271) );
  OR3_X1 U39 ( .A1(B[14]), .A2(B[15]), .A3(n267), .ZN(n265) );
  NAND2_X1 U40 ( .A1(n202), .A2(n293), .ZN(n241) );
  NOR3_X1 U41 ( .A1(B[36]), .A2(B[37]), .A3(n244), .ZN(n202) );
  INV_X1 U42 ( .A(n248), .ZN(n296) );
  XNOR2_X1 U43 ( .A(B[37]), .B(n245), .ZN(DIFF[37]) );
  NOR2_X1 U44 ( .A1(B[36]), .A2(n244), .ZN(n245) );
  XNOR2_X1 U45 ( .A(n262), .B(B[33]), .ZN(DIFF[33]) );
  NOR2_X1 U46 ( .A1(n248), .A2(B[32]), .ZN(n262) );
  NOR3_X1 U47 ( .A1(B[36]), .A2(B[37]), .A3(n244), .ZN(n243) );
  OR3_X1 U48 ( .A1(B[32]), .A2(B[33]), .A3(n248), .ZN(n247) );
  XNOR2_X1 U49 ( .A(n228), .B(B[45]), .ZN(DIFF[45]) );
  NOR2_X1 U50 ( .A1(n235), .A2(B[44]), .ZN(n228) );
  XNOR2_X1 U51 ( .A(n254), .B(B[29]), .ZN(DIFF[29]) );
  NOR2_X1 U52 ( .A1(n252), .A2(B[28]), .ZN(n254) );
  XNOR2_X1 U53 ( .A(n241), .B(n294), .ZN(DIFF[39]) );
  XNOR2_X1 U54 ( .A(n213), .B(B[49]), .ZN(DIFF[49]) );
  NOR2_X1 U55 ( .A1(n231), .A2(B[48]), .ZN(n213) );
  XNOR2_X1 U56 ( .A(B[47]), .B(n234), .ZN(DIFF[47]) );
  NOR2_X1 U57 ( .A1(B[46]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U58 ( .A(B[31]), .B(n251), .ZN(DIFF[31]) );
  NOR2_X1 U59 ( .A1(B[30]), .A2(n250), .ZN(n251) );
  XNOR2_X1 U64 ( .A(n224), .B(B[57]), .ZN(DIFF[57]) );
  NOR2_X1 U65 ( .A1(n223), .A2(B[56]), .ZN(n224) );
  XNOR2_X1 U66 ( .A(B[55]), .B(n226), .ZN(DIFF[55]) );
  NOR2_X1 U67 ( .A1(B[54]), .A2(n225), .ZN(n226) );
  XNOR2_X1 U68 ( .A(n219), .B(B[53]), .ZN(DIFF[53]) );
  NOR2_X1 U69 ( .A1(n227), .A2(B[52]), .ZN(n219) );
  XNOR2_X1 U70 ( .A(B[51]), .B(n230), .ZN(DIFF[51]) );
  NOR2_X1 U71 ( .A1(B[50]), .A2(n229), .ZN(n230) );
  XNOR2_X1 U72 ( .A(B[27]), .B(n256), .ZN(DIFF[27]) );
  NOR2_X1 U73 ( .A1(B[26]), .A2(n255), .ZN(n256) );
  XNOR2_X1 U74 ( .A(n240), .B(B[25]), .ZN(DIFF[25]) );
  NOR2_X1 U75 ( .A1(n257), .A2(B[24]), .ZN(n240) );
  XNOR2_X1 U76 ( .A(n258), .B(B[21]), .ZN(DIFF[21]) );
  NOR2_X1 U77 ( .A1(n261), .A2(B[20]), .ZN(n258) );
  XNOR2_X1 U78 ( .A(B[59]), .B(n222), .ZN(DIFF[59]) );
  NOR2_X1 U79 ( .A1(B[58]), .A2(n220), .ZN(n222) );
  XNOR2_X1 U80 ( .A(B[23]), .B(n260), .ZN(DIFF[23]) );
  NOR2_X1 U81 ( .A1(B[22]), .A2(n259), .ZN(n260) );
  XNOR2_X1 U82 ( .A(B[17]), .B(n266), .ZN(DIFF[17]) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(n265), .ZN(n266) );
  XNOR2_X1 U84 ( .A(n236), .B(B[61]), .ZN(DIFF[61]) );
  NOR2_X1 U85 ( .A1(n218), .A2(B[60]), .ZN(n236) );
  NAND2_X1 U86 ( .A1(n217), .A2(n295), .ZN(n216) );
  XNOR2_X1 U87 ( .A(B[43]), .B(n238), .ZN(DIFF[43]) );
  NOR2_X1 U88 ( .A1(B[42]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U89 ( .A(n232), .B(B[41]), .ZN(DIFF[41]) );
  NOR2_X1 U90 ( .A1(n239), .A2(B[40]), .ZN(n232) );
  NOR3_X1 U91 ( .A1(n221), .A2(B[4]), .A3(n284), .ZN(n212) );
  OR3_X1 U92 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n284) );
  XNOR2_X1 U93 ( .A(n268), .B(B[7]), .ZN(DIFF[7]) );
  NOR2_X1 U94 ( .A1(n214), .A2(B[6]), .ZN(n268) );
  NOR2_X1 U95 ( .A1(n221), .A2(B[4]), .ZN(n215) );
  XNOR2_X1 U96 ( .A(n215), .B(B[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U99 ( .A(n253), .B(B[2]), .ZN(DIFF[2]) );
  OR2_X1 U102 ( .A1(n242), .A2(B[3]), .ZN(n221) );
  NAND2_X1 U105 ( .A1(n215), .A2(n299), .ZN(n214) );
  INV_X1 U109 ( .A(B[5]), .ZN(n299) );
  NAND2_X1 U112 ( .A1(n253), .A2(n298), .ZN(n242) );
  INV_X1 U115 ( .A(B[2]), .ZN(n298) );
  NOR2_X1 U118 ( .A1(B[1]), .A2(B[0]), .ZN(n253) );
  INV_X1 U121 ( .A(B[9]), .ZN(n285) );
  INV_X1 U124 ( .A(B[10]), .ZN(n286) );
  INV_X1 U127 ( .A(B[12]), .ZN(n287) );
  INV_X1 U130 ( .A(B[18]), .ZN(n288) );
  INV_X1 U135 ( .A(B[32]), .ZN(n289) );
  INV_X1 U140 ( .A(B[33]), .ZN(n290) );
  INV_X1 U141 ( .A(B[34]), .ZN(n291) );
  INV_X1 U142 ( .A(B[35]), .ZN(n292) );
  INV_X1 U143 ( .A(B[38]), .ZN(n293) );
  INV_X1 U144 ( .A(B[39]), .ZN(n294) );
  INV_X1 U145 ( .A(B[62]), .ZN(n295) );
endmodule


module complement_NBIT64_25 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_25_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_24_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n215, n216, n217, n219, n220, n221, n223, n224, n225, n227,
         n228, n229, n231, n232, n233, n234, n235, n236, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n253, n254, n255, n256, n257, n259, n260, n261, n262, n263, n264,
         n265, n266, n194, n195, n196, n197, n198, n199, n200, n201, n268,
         n269, n270, n271, n272, n273, n274, n275, n276;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U96 ( .A(n204), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U97 ( .A(n206), .B(B[6]), .Z(DIFF[6]) );
  NAND3_X1 U98 ( .A1(n275), .A2(n276), .A3(n207), .ZN(n206) );
  XOR2_X1 U99 ( .A(n208), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U100 ( .A(n210), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U101 ( .A(n213), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U103 ( .A(n212), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U104 ( .A(n215), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U106 ( .A(n217), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U107 ( .A(n219), .B(B[52]), .Z(DIFF[52]) );
  XOR2_X1 U109 ( .A(n221), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U110 ( .A(n223), .B(B[48]), .Z(DIFF[48]) );
  XOR2_X1 U112 ( .A(n225), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U113 ( .A(n227), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U115 ( .A(n229), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U116 ( .A(n231), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U117 ( .A(n234), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U118 ( .A(n235), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U120 ( .A(n236), .B(B[36]), .Z(DIFF[36]) );
  XOR2_X1 U121 ( .A(n238), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U122 ( .A(n240), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U123 ( .A(n243), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U124 ( .A(n242), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U125 ( .A(n244), .B(B[28]), .Z(DIFF[28]) );
  XOR2_X1 U126 ( .A(n248), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U127 ( .A(n247), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U128 ( .A(n249), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U130 ( .A(n251), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U131 ( .A(n253), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U132 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U133 ( .A(n256), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U135 ( .A(n257), .B(B[16]), .Z(DIFF[16]) );
  XOR2_X1 U136 ( .A(n259), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U137 ( .A(n265), .B(B[10]), .Z(DIFF[10]) );
  NAND3_X1 U138 ( .A1(n207), .A2(n275), .A3(n266), .ZN(n204) );
  XOR2_X1 U4 ( .A(n209), .B(n273), .Z(DIFF[62]) );
  XOR2_X1 U39 ( .A(n272), .B(n233), .Z(DIFF[39]) );
  XOR2_X1 U45 ( .A(n270), .B(n255), .Z(DIFF[19]) );
  XOR2_X1 U47 ( .A(n239), .B(n271), .Z(DIFF[34]) );
  XOR2_X1 U48 ( .A(n269), .B(n261), .Z(DIFF[13]) );
  OR3_X1 U3 ( .A1(B[44]), .A2(B[45]), .A3(n227), .ZN(n225) );
  OR3_X1 U5 ( .A1(B[36]), .A2(B[37]), .A3(n236), .ZN(n235) );
  OR3_X1 U6 ( .A1(B[30]), .A2(B[31]), .A3(n242), .ZN(n240) );
  NOR3_X1 U7 ( .A1(B[60]), .A2(B[61]), .A3(n210), .ZN(n209) );
  OR3_X1 U8 ( .A1(B[58]), .A2(B[59]), .A3(n212), .ZN(n210) );
  OR3_X1 U9 ( .A1(B[42]), .A2(B[43]), .A3(n229), .ZN(n227) );
  OR3_X1 U10 ( .A1(B[46]), .A2(B[47]), .A3(n225), .ZN(n223) );
  OR3_X1 U11 ( .A1(B[50]), .A2(B[51]), .A3(n221), .ZN(n219) );
  OR3_X1 U12 ( .A1(B[54]), .A2(B[55]), .A3(n217), .ZN(n215) );
  OR3_X1 U13 ( .A1(B[48]), .A2(B[49]), .A3(n223), .ZN(n221) );
  OR3_X1 U14 ( .A1(B[52]), .A2(B[53]), .A3(n219), .ZN(n217) );
  OR3_X1 U15 ( .A1(B[56]), .A2(B[57]), .A3(n215), .ZN(n212) );
  OR3_X1 U16 ( .A1(B[40]), .A2(B[41]), .A3(n231), .ZN(n229) );
  XNOR2_X1 U17 ( .A(B[9]), .B(n203), .ZN(DIFF[9]) );
  NAND2_X1 U18 ( .A1(n261), .A2(n269), .ZN(n259) );
  NAND2_X1 U19 ( .A1(n233), .A2(n272), .ZN(n231) );
  NAND2_X1 U20 ( .A1(n255), .A2(n270), .ZN(n253) );
  NAND2_X1 U21 ( .A1(n239), .A2(n271), .ZN(n238) );
  NAND2_X1 U22 ( .A1(n203), .A2(n268), .ZN(n265) );
  OR3_X1 U23 ( .A1(B[28]), .A2(B[29]), .A3(n244), .ZN(n242) );
  NOR3_X1 U24 ( .A1(n204), .A2(B[12]), .A3(n262), .ZN(n261) );
  NOR3_X1 U25 ( .A1(B[32]), .A2(B[33]), .A3(n240), .ZN(n239) );
  NOR2_X1 U26 ( .A1(n204), .A2(B[8]), .ZN(n203) );
  NOR2_X1 U27 ( .A1(n256), .A2(B[18]), .ZN(n255) );
  NOR2_X1 U28 ( .A1(n235), .A2(B[38]), .ZN(n233) );
  XNOR2_X1 U29 ( .A(B[12]), .B(n263), .ZN(DIFF[12]) );
  NOR2_X1 U30 ( .A1(n204), .A2(n262), .ZN(n263) );
  XNOR2_X1 U31 ( .A(B[15]), .B(n260), .ZN(DIFF[15]) );
  NOR2_X1 U32 ( .A1(B[14]), .A2(n259), .ZN(n260) );
  OR4_X1 U33 ( .A1(B[10]), .A2(B[11]), .A3(B[8]), .A4(B[9]), .ZN(n262) );
  OR2_X1 U34 ( .A1(n238), .A2(B[35]), .ZN(n236) );
  OR3_X1 U35 ( .A1(B[22]), .A2(B[23]), .A3(n251), .ZN(n249) );
  OR3_X1 U36 ( .A1(B[26]), .A2(B[27]), .A3(n247), .ZN(n244) );
  OR3_X1 U37 ( .A1(B[20]), .A2(B[21]), .A3(n253), .ZN(n251) );
  OR3_X1 U38 ( .A1(B[14]), .A2(B[15]), .A3(n259), .ZN(n257) );
  OR3_X1 U40 ( .A1(B[24]), .A2(B[25]), .A3(n249), .ZN(n247) );
  OR3_X1 U41 ( .A1(B[16]), .A2(B[17]), .A3(n257), .ZN(n256) );
  XNOR2_X1 U42 ( .A(n199), .B(B[37]), .ZN(DIFF[37]) );
  NOR2_X1 U43 ( .A1(n236), .A2(B[36]), .ZN(n199) );
  XNOR2_X1 U44 ( .A(B[53]), .B(n220), .ZN(DIFF[53]) );
  NOR2_X1 U46 ( .A1(B[52]), .A2(n219), .ZN(n220) );
  XNOR2_X1 U49 ( .A(n195), .B(B[55]), .ZN(DIFF[55]) );
  NOR2_X1 U50 ( .A1(n217), .A2(B[54]), .ZN(n195) );
  XNOR2_X1 U51 ( .A(B[49]), .B(n224), .ZN(DIFF[49]) );
  NOR2_X1 U52 ( .A1(B[48]), .A2(n223), .ZN(n224) );
  XNOR2_X1 U53 ( .A(B[45]), .B(n228), .ZN(DIFF[45]) );
  NOR2_X1 U54 ( .A1(B[44]), .A2(n227), .ZN(n228) );
  XNOR2_X1 U55 ( .A(n194), .B(B[51]), .ZN(DIFF[51]) );
  NOR2_X1 U56 ( .A1(n221), .A2(B[50]), .ZN(n194) );
  XNOR2_X1 U57 ( .A(B[57]), .B(n216), .ZN(DIFF[57]) );
  NOR2_X1 U58 ( .A1(B[56]), .A2(n215), .ZN(n216) );
  OR2_X1 U59 ( .A1(n247), .A2(B[26]), .ZN(n248) );
  XNOR2_X1 U60 ( .A(n200), .B(B[23]), .ZN(DIFF[23]) );
  NOR2_X1 U61 ( .A1(n251), .A2(B[22]), .ZN(n200) );
  XNOR2_X1 U62 ( .A(B[11]), .B(n264), .ZN(DIFF[11]) );
  NOR2_X1 U63 ( .A1(B[10]), .A2(n265), .ZN(n264) );
  XNOR2_X1 U64 ( .A(n198), .B(B[43]), .ZN(DIFF[43]) );
  NOR2_X1 U65 ( .A1(n229), .A2(B[42]), .ZN(n198) );
  OR2_X1 U66 ( .A1(n242), .A2(B[30]), .ZN(n243) );
  XNOR2_X1 U67 ( .A(B[33]), .B(n241), .ZN(DIFF[33]) );
  NOR2_X1 U68 ( .A1(B[32]), .A2(n240), .ZN(n241) );
  XNOR2_X1 U69 ( .A(n196), .B(B[59]), .ZN(DIFF[59]) );
  NOR2_X1 U70 ( .A1(n212), .A2(B[58]), .ZN(n196) );
  XNOR2_X1 U71 ( .A(B[41]), .B(n232), .ZN(DIFF[41]) );
  NOR2_X1 U72 ( .A1(B[40]), .A2(n231), .ZN(n232) );
  XNOR2_X1 U73 ( .A(n197), .B(B[47]), .ZN(DIFF[47]) );
  NOR2_X1 U74 ( .A1(n225), .A2(B[46]), .ZN(n197) );
  XNOR2_X1 U75 ( .A(B[21]), .B(n254), .ZN(DIFF[21]) );
  NOR2_X1 U76 ( .A1(B[20]), .A2(n253), .ZN(n254) );
  XNOR2_X1 U77 ( .A(B[29]), .B(n246), .ZN(DIFF[29]) );
  NOR2_X1 U78 ( .A1(B[28]), .A2(n244), .ZN(n246) );
  XNOR2_X1 U79 ( .A(n201), .B(B[17]), .ZN(DIFF[17]) );
  NOR2_X1 U80 ( .A1(n257), .A2(B[16]), .ZN(n201) );
  XNOR2_X1 U81 ( .A(B[61]), .B(n211), .ZN(DIFF[61]) );
  NOR2_X1 U82 ( .A1(B[60]), .A2(n210), .ZN(n211) );
  NAND2_X1 U83 ( .A1(n209), .A2(n273), .ZN(n208) );
  XNOR2_X1 U84 ( .A(B[25]), .B(n250), .ZN(DIFF[25]) );
  NOR2_X1 U85 ( .A1(B[24]), .A2(n249), .ZN(n250) );
  NOR3_X1 U86 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n266) );
  NOR2_X1 U87 ( .A1(n234), .A2(B[3]), .ZN(n207) );
  NAND2_X1 U88 ( .A1(n207), .A2(n275), .ZN(n213) );
  INV_X1 U89 ( .A(B[5]), .ZN(n276) );
  XNOR2_X1 U90 ( .A(B[7]), .B(n205), .ZN(DIFF[7]) );
  NOR2_X1 U91 ( .A1(B[6]), .A2(n206), .ZN(n205) );
  XNOR2_X1 U92 ( .A(n245), .B(B[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U93 ( .A(n207), .B(B[4]), .ZN(DIFF[4]) );
  NAND2_X1 U94 ( .A1(n245), .A2(n274), .ZN(n234) );
  INV_X1 U95 ( .A(B[2]), .ZN(n274) );
  INV_X1 U102 ( .A(B[4]), .ZN(n275) );
  NOR2_X1 U105 ( .A1(B[1]), .A2(\B[0] ), .ZN(n245) );
  INV_X1 U108 ( .A(B[9]), .ZN(n268) );
  INV_X1 U111 ( .A(B[13]), .ZN(n269) );
  INV_X1 U114 ( .A(B[19]), .ZN(n270) );
  INV_X1 U119 ( .A(B[34]), .ZN(n271) );
  INV_X1 U129 ( .A(B[39]), .ZN(n272) );
  INV_X1 U134 ( .A(B[62]), .ZN(n273) );
endmodule


module complement_NBIT64_24 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_24_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_23_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n9, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n50, n52, n55, n56, n58, n60, n62, n63, n68, n71,
         n74, n75, n80, n83, n86, n87, n92, n96, n99, n100, n102, n103, n104,
         n108, n110, n111, n113, n115, n120, n121, n131, n132, n134, n135,
         n136, n137, n140, n141, n142, n145, n146, n148, n149, n150, n152,
         n154, n155, n160, n162, n165, n166, n173, n174, n175, n177, n178,
         n179, n183, n184, n187, n188, n189, n193, n195, n196, n201, n202,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U9 ( .A(n4), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U11 ( .A(n5), .B(n299), .Z(DIFF[12]) );
  XOR2_X1 U13 ( .A(n365), .B(n6), .Z(DIFF[3]) );
  XOR2_X1 U15 ( .A(n7), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U37 ( .A(n9), .B(n328), .Z(DIFF[41]) );
  XOR2_X1 U38 ( .A(B[43]), .B(n120), .Z(DIFF[43]) );
  XOR2_X1 U47 ( .A(n92), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U52 ( .A(n346), .B(n356), .Z(DIFF[57]) );
  XOR2_X1 U53 ( .A(n342), .B(n355), .Z(DIFF[53]) );
  XOR2_X1 U58 ( .A(n338), .B(n354), .Z(DIFF[49]) );
  XOR2_X1 U59 ( .A(n113), .B(n332), .Z(DIFF[44]) );
  XOR2_X1 U60 ( .A(n80), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U64 ( .A(n68), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U85 ( .A(n162), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U89 ( .A(n11), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U94 ( .A(n1), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U95 ( .A(n175), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U96 ( .A(B[40]), .B(n115), .Z(DIFF[40]) );
  XOR2_X1 U116 ( .A(B[31]), .B(n154), .Z(DIFF[31]) );
  XOR2_X1 U121 ( .A(n307), .B(n352), .Z(DIFF[20]) );
  XOR2_X1 U151 ( .A(B[15]), .B(n193), .Z(DIFF[15]) );
  XOR2_X1 U155 ( .A(B[19]), .B(n183), .Z(DIFF[19]) );
  XOR2_X1 U164 ( .A(B[10]), .B(n205), .Z(DIFF[10]) );
  XOR2_X1 U167 ( .A(B[14]), .B(n196), .Z(DIFF[14]) );
  XOR2_X1 U169 ( .A(B[27]), .B(n165), .Z(DIFF[27]) );
  XOR2_X1 U175 ( .A(B[23]), .B(n173), .Z(DIFF[23]) );
  XOR2_X1 U177 ( .A(B[35]), .B(n140), .Z(DIFF[35]) );
  XOR2_X1 U179 ( .A(B[39]), .B(n131), .Z(DIFF[39]) );
  XOR2_X1 U181 ( .A(B[9]), .B(n50), .Z(DIFF[9]) );
  XOR2_X1 U189 ( .A(n364), .B(n19), .Z(DIFF[2]) );
  XOR2_X1 U190 ( .A(n18), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U191 ( .A(n52), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U192 ( .A(n368), .B(n2), .Z(DIFF[8]) );
  XOR2_X1 U193 ( .A(n367), .B(n55), .Z(DIFF[6]) );
  XOR2_X1 U200 ( .A(\B[0] ), .B(B[1]), .Z(DIFF[1]) );
  NAND3_X1 U247 ( .A1(n368), .A2(n20), .A3(n361), .ZN(n50) );
  NAND3_X1 U248 ( .A1(n347), .A2(n348), .A3(n346), .ZN(n63) );
  NAND3_X1 U250 ( .A1(n343), .A2(n344), .A3(n342), .ZN(n75) );
  NAND3_X1 U252 ( .A1(n339), .A2(n340), .A3(n338), .ZN(n87) );
  NAND3_X1 U254 ( .A1(n359), .A2(n17), .A3(n102), .ZN(n100) );
  NAND3_X1 U261 ( .A1(n358), .A2(n16), .A3(n148), .ZN(n146) );
  NAND3_X1 U267 ( .A1(n301), .A2(n302), .A3(n357), .ZN(n193) );
  NAND3_X1 U268 ( .A1(n2), .A2(n301), .A3(n14), .ZN(n196) );
  XOR2_X1 U3 ( .A(n208), .B(n344), .Z(DIFF[55]) );
  XOR2_X1 U5 ( .A(n209), .B(n348), .Z(DIFF[59]) );
  XOR2_X1 U7 ( .A(n210), .B(n340), .Z(DIFF[51]) );
  XOR2_X1 U32 ( .A(n83), .B(n341), .Z(DIFF[52]) );
  XOR2_X1 U33 ( .A(n71), .B(n345), .Z(DIFF[56]) );
  XOR2_X1 U36 ( .A(n349), .B(n60), .Z(DIFF[60]) );
  XOR2_X1 U39 ( .A(n56), .B(n351), .Z(DIFF[62]) );
  XOR2_X1 U40 ( .A(n350), .B(n58), .Z(DIFF[61]) );
  XOR2_X1 U50 ( .A(n96), .B(n337), .Z(DIFF[48]) );
  XOR2_X1 U51 ( .A(n211), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U91 ( .A(n3), .B(n303), .Z(DIFF[16]) );
  XOR2_X1 U92 ( .A(n353), .B(n323), .Z(DIFF[36]) );
  INV_X1 U4 ( .A(n74), .ZN(n355) );
  INV_X1 U6 ( .A(n62), .ZN(n356) );
  NAND2_X1 U8 ( .A1(n83), .A2(n341), .ZN(n74) );
  NOR2_X1 U10 ( .A1(n92), .A2(B[50]), .ZN(n210) );
  NOR2_X1 U12 ( .A1(n80), .A2(B[54]), .ZN(n208) );
  AND2_X1 U14 ( .A1(n111), .A2(n334), .ZN(n110) );
  NAND2_X1 U16 ( .A1(n338), .A2(n354), .ZN(n92) );
  NAND2_X1 U17 ( .A1(n342), .A2(n355), .ZN(n80) );
  NAND2_X1 U18 ( .A1(n333), .A2(n334), .ZN(n104) );
  NOR2_X1 U19 ( .A1(n74), .A2(n75), .ZN(n71) );
  NOR2_X1 U20 ( .A1(n62), .A2(n63), .ZN(n60) );
  NAND2_X1 U21 ( .A1(n71), .A2(n345), .ZN(n62) );
  NOR2_X1 U22 ( .A1(n68), .A2(B[58]), .ZN(n209) );
  NAND2_X1 U23 ( .A1(n346), .A2(n356), .ZN(n68) );
  AND2_X1 U24 ( .A1(n350), .A2(n58), .ZN(n56) );
  AND2_X1 U25 ( .A1(n349), .A2(n60), .ZN(n58) );
  NOR2_X1 U26 ( .A1(n1), .A2(B[29]), .ZN(n155) );
  NOR2_X1 U27 ( .A1(n9), .A2(n328), .ZN(n121) );
  NOR2_X1 U28 ( .A1(n113), .A2(n332), .ZN(n111) );
  NOR2_X1 U29 ( .A1(n86), .A2(n87), .ZN(n83) );
  NAND4_X1 U30 ( .A1(n327), .A2(n331), .A3(n330), .A4(n329), .ZN(n108) );
  XNOR2_X1 U31 ( .A(B[45]), .B(n111), .ZN(DIFF[45]) );
  XNOR2_X1 U34 ( .A(n121), .B(B[42]), .ZN(DIFF[42]) );
  XNOR2_X1 U35 ( .A(n110), .B(B[46]), .ZN(DIFF[46]) );
  INV_X1 U41 ( .A(n86), .ZN(n354) );
  NAND2_X1 U42 ( .A1(n335), .A2(n336), .ZN(n103) );
  NAND2_X1 U43 ( .A1(n330), .A2(n121), .ZN(n120) );
  NAND2_X1 U44 ( .A1(n335), .A2(n110), .ZN(n4) );
  NAND2_X1 U45 ( .A1(n56), .A2(n351), .ZN(n211) );
  NOR2_X1 U46 ( .A1(n175), .A2(B[21]), .ZN(n174) );
  NOR2_X1 U48 ( .A1(n11), .A2(B[25]), .ZN(n166) );
  XNOR2_X1 U49 ( .A(n301), .B(n195), .ZN(DIFF[13]) );
  INV_X1 U54 ( .A(n145), .ZN(n352) );
  AND2_X1 U55 ( .A1(n142), .A2(n320), .ZN(n141) );
  NAND2_X1 U56 ( .A1(n160), .A2(n315), .ZN(n1) );
  NAND2_X1 U57 ( .A1(n352), .A2(n307), .ZN(n175) );
  OR2_X1 U61 ( .A1(B[24]), .A2(n162), .ZN(n11) );
  NAND2_X1 U62 ( .A1(n315), .A2(n316), .ZN(n150) );
  NAND2_X1 U63 ( .A1(n96), .A2(n337), .ZN(n86) );
  INV_X1 U65 ( .A(n99), .ZN(n353) );
  OR2_X1 U66 ( .A1(B[40]), .A2(n115), .ZN(n9) );
  OR2_X1 U67 ( .A1(n108), .A2(n115), .ZN(n113) );
  NOR2_X1 U68 ( .A1(n145), .A2(n146), .ZN(n134) );
  NOR2_X1 U69 ( .A1(n149), .A2(n150), .ZN(n148) );
  INV_X1 U70 ( .A(n152), .ZN(n358) );
  NAND2_X1 U71 ( .A1(n15), .A2(n2), .ZN(n5) );
  NOR2_X1 U72 ( .A1(n162), .A2(n152), .ZN(n160) );
  XNOR2_X1 U73 ( .A(B[28]), .B(n160), .ZN(DIFF[28]) );
  XNOR2_X1 U74 ( .A(n155), .B(B[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U75 ( .A(n166), .B(B[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U76 ( .A(B[33]), .B(n142), .ZN(DIFF[33]) );
  XNOR2_X1 U77 ( .A(n212), .B(n298), .ZN(DIFF[11]) );
  NAND2_X1 U78 ( .A1(n201), .A2(n202), .ZN(n212) );
  NOR2_X1 U79 ( .A1(n366), .A2(B[10]), .ZN(n202) );
  NOR2_X1 U80 ( .A1(n204), .A2(n52), .ZN(n201) );
  NAND2_X1 U81 ( .A1(n16), .A2(n352), .ZN(n162) );
  NAND2_X1 U82 ( .A1(n14), .A2(n2), .ZN(n195) );
  NAND2_X1 U83 ( .A1(n3), .A2(n177), .ZN(n145) );
  NOR2_X1 U84 ( .A1(n178), .A2(n179), .ZN(n177) );
  NAND2_X1 U86 ( .A1(n303), .A2(n306), .ZN(n178) );
  NAND2_X1 U87 ( .A1(n304), .A2(n305), .ZN(n179) );
  AND2_X1 U88 ( .A1(n13), .A2(n304), .ZN(n184) );
  AND2_X1 U90 ( .A1(n319), .A2(n134), .ZN(n142) );
  AND2_X1 U93 ( .A1(n3), .A2(n303), .ZN(n13) );
  AND2_X1 U97 ( .A1(n15), .A2(n300), .ZN(n14) );
  NOR2_X1 U98 ( .A1(n99), .A2(n100), .ZN(n96) );
  NOR2_X1 U99 ( .A1(n103), .A2(n104), .ZN(n102) );
  INV_X1 U100 ( .A(n108), .ZN(n359) );
  XNOR2_X1 U101 ( .A(n132), .B(B[38]), .ZN(DIFF[38]) );
  NAND2_X1 U102 ( .A1(n134), .A2(n135), .ZN(n99) );
  NOR2_X1 U103 ( .A1(n136), .A2(n137), .ZN(n135) );
  NAND2_X1 U104 ( .A1(n319), .A2(n322), .ZN(n136) );
  NAND2_X1 U105 ( .A1(n320), .A2(n321), .ZN(n137) );
  AND2_X1 U106 ( .A1(n12), .A2(n324), .ZN(n132) );
  NAND2_X1 U107 ( .A1(n17), .A2(n353), .ZN(n115) );
  AND2_X1 U108 ( .A1(n353), .A2(n323), .ZN(n12) );
  INV_X1 U109 ( .A(n52), .ZN(n361) );
  NAND2_X1 U110 ( .A1(n305), .A2(n184), .ZN(n183) );
  NAND2_X1 U111 ( .A1(n309), .A2(n174), .ZN(n173) );
  NAND2_X1 U112 ( .A1(n317), .A2(n155), .ZN(n154) );
  NAND2_X1 U113 ( .A1(n321), .A2(n141), .ZN(n140) );
  NAND4_X1 U114 ( .A1(n311), .A2(n314), .A3(n313), .A4(n312), .ZN(n152) );
  XNOR2_X1 U115 ( .A(B[17]), .B(n13), .ZN(DIFF[17]) );
  XNOR2_X1 U117 ( .A(n174), .B(B[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U118 ( .A(B[32]), .B(n134), .ZN(DIFF[32]) );
  XNOR2_X1 U119 ( .A(n184), .B(B[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U120 ( .A(n141), .B(B[34]), .ZN(DIFF[34]) );
  AND3_X1 U122 ( .A1(n187), .A2(n188), .A3(n15), .ZN(n3) );
  NOR2_X1 U123 ( .A1(n299), .A2(n52), .ZN(n187) );
  NOR3_X1 U124 ( .A1(n189), .A2(n366), .A3(B[15]), .ZN(n188) );
  NAND2_X1 U125 ( .A1(n301), .A2(n302), .ZN(n189) );
  NAND2_X1 U126 ( .A1(n368), .A2(n296), .ZN(n204) );
  AND4_X1 U127 ( .A1(n298), .A2(n297), .A3(n296), .A4(n368), .ZN(n15) );
  AND4_X1 U128 ( .A1(n307), .A2(n310), .A3(n309), .A4(n308), .ZN(n16) );
  NAND2_X1 U129 ( .A1(n317), .A2(n318), .ZN(n149) );
  NAND2_X1 U130 ( .A1(n313), .A2(n166), .ZN(n165) );
  NAND2_X1 U131 ( .A1(n325), .A2(n132), .ZN(n131) );
  XNOR2_X1 U132 ( .A(B[37]), .B(n12), .ZN(DIFF[37]) );
  AND4_X1 U133 ( .A1(n323), .A2(n326), .A3(n325), .A4(n324), .ZN(n17) );
  AND2_X1 U134 ( .A1(n361), .A2(n20), .ZN(n2) );
  INV_X1 U135 ( .A(n20), .ZN(n366) );
  NAND4_X1 U136 ( .A1(n363), .A2(n362), .A3(n364), .A4(n365), .ZN(n52) );
  AND2_X1 U137 ( .A1(n363), .A2(n362), .ZN(n19) );
  NAND4_X1 U138 ( .A1(n206), .A2(n20), .A3(n207), .A4(n365), .ZN(n205) );
  NOR2_X1 U139 ( .A1(B[1]), .A2(B[2]), .ZN(n207) );
  NOR2_X1 U140 ( .A1(n204), .A2(\B[0] ), .ZN(n206) );
  INV_X1 U141 ( .A(n195), .ZN(n357) );
  NOR2_X1 U142 ( .A1(n18), .A2(B[5]), .ZN(n55) );
  NAND2_X1 U143 ( .A1(n367), .A2(n55), .ZN(n7) );
  NOR2_X1 U144 ( .A1(n360), .A2(B[2]), .ZN(n6) );
  INV_X1 U145 ( .A(n19), .ZN(n360) );
  AND2_X1 U146 ( .A1(n213), .A2(n214), .ZN(n20) );
  NOR2_X1 U147 ( .A1(B[5]), .A2(B[4]), .ZN(n213) );
  NOR2_X1 U148 ( .A1(B[7]), .A2(B[6]), .ZN(n214) );
  OR2_X1 U149 ( .A1(B[4]), .A2(n52), .ZN(n18) );
  INV_X1 U150 ( .A(B[8]), .ZN(n368) );
  INV_X1 U152 ( .A(B[3]), .ZN(n365) );
  INV_X1 U153 ( .A(B[2]), .ZN(n364) );
  INV_X1 U154 ( .A(B[6]), .ZN(n367) );
  INV_X1 U156 ( .A(\B[0] ), .ZN(n362) );
  INV_X1 U157 ( .A(B[1]), .ZN(n363) );
  INV_X1 U158 ( .A(B[9]), .ZN(n296) );
  INV_X1 U159 ( .A(B[10]), .ZN(n297) );
  INV_X1 U160 ( .A(B[11]), .ZN(n298) );
  INV_X1 U161 ( .A(n300), .ZN(n299) );
  INV_X1 U162 ( .A(B[12]), .ZN(n300) );
  INV_X1 U163 ( .A(B[13]), .ZN(n301) );
  INV_X1 U165 ( .A(B[14]), .ZN(n302) );
  INV_X1 U166 ( .A(B[16]), .ZN(n303) );
  INV_X1 U168 ( .A(B[17]), .ZN(n304) );
  INV_X1 U170 ( .A(B[18]), .ZN(n305) );
  INV_X1 U171 ( .A(B[19]), .ZN(n306) );
  INV_X1 U172 ( .A(B[20]), .ZN(n307) );
  INV_X1 U173 ( .A(B[21]), .ZN(n308) );
  INV_X1 U174 ( .A(B[22]), .ZN(n309) );
  INV_X1 U176 ( .A(B[23]), .ZN(n310) );
  INV_X1 U178 ( .A(B[24]), .ZN(n311) );
  INV_X1 U180 ( .A(B[25]), .ZN(n312) );
  INV_X1 U182 ( .A(B[26]), .ZN(n313) );
  INV_X1 U183 ( .A(B[27]), .ZN(n314) );
  INV_X1 U184 ( .A(B[28]), .ZN(n315) );
  INV_X1 U185 ( .A(B[29]), .ZN(n316) );
  INV_X1 U186 ( .A(B[30]), .ZN(n317) );
  INV_X1 U187 ( .A(B[31]), .ZN(n318) );
  INV_X1 U188 ( .A(B[32]), .ZN(n319) );
  INV_X1 U194 ( .A(B[33]), .ZN(n320) );
  INV_X1 U195 ( .A(B[34]), .ZN(n321) );
  INV_X1 U196 ( .A(B[35]), .ZN(n322) );
  INV_X1 U197 ( .A(B[36]), .ZN(n323) );
  INV_X1 U198 ( .A(B[37]), .ZN(n324) );
  INV_X1 U199 ( .A(B[38]), .ZN(n325) );
  INV_X1 U201 ( .A(B[39]), .ZN(n326) );
  INV_X1 U202 ( .A(B[40]), .ZN(n327) );
  INV_X1 U203 ( .A(n329), .ZN(n328) );
  INV_X1 U204 ( .A(B[41]), .ZN(n329) );
  INV_X1 U205 ( .A(B[42]), .ZN(n330) );
  INV_X1 U206 ( .A(B[43]), .ZN(n331) );
  INV_X1 U207 ( .A(n333), .ZN(n332) );
  INV_X1 U208 ( .A(B[44]), .ZN(n333) );
  INV_X1 U209 ( .A(B[45]), .ZN(n334) );
  INV_X1 U210 ( .A(B[46]), .ZN(n335) );
  INV_X1 U211 ( .A(B[47]), .ZN(n336) );
  INV_X1 U212 ( .A(B[48]), .ZN(n337) );
  INV_X1 U213 ( .A(B[49]), .ZN(n338) );
  INV_X1 U214 ( .A(B[50]), .ZN(n339) );
  INV_X1 U215 ( .A(B[51]), .ZN(n340) );
  INV_X1 U216 ( .A(B[52]), .ZN(n341) );
  INV_X1 U217 ( .A(B[53]), .ZN(n342) );
  INV_X1 U218 ( .A(B[54]), .ZN(n343) );
  INV_X1 U219 ( .A(B[55]), .ZN(n344) );
  INV_X1 U220 ( .A(B[56]), .ZN(n345) );
  INV_X1 U221 ( .A(B[57]), .ZN(n346) );
  INV_X1 U222 ( .A(B[58]), .ZN(n347) );
  INV_X1 U223 ( .A(B[59]), .ZN(n348) );
  INV_X1 U224 ( .A(B[60]), .ZN(n349) );
  INV_X1 U225 ( .A(B[61]), .ZN(n350) );
  INV_X1 U226 ( .A(B[62]), .ZN(n351) );
endmodule


module complement_NBIT64_23 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_23_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_22_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15,
         n16, n19, n20, n21, n22, n24, n25, n26, n27, n28, n36, n39, n40, n43,
         n45, n47, n48, n53, n55, n57, n58, n62, n64, n66, n67, n71, n73, n74,
         n76, n77, n79, n80, n81, n86, n88, n92, n98, n107, n111, n112, n114,
         n115, n116, n117, n123, n124, n127, n128, n130, n131, n132, n137,
         n138, n139, n140, n143, n149, n150, n151, n158, n159, n160, n162,
         n163, n164, n165, n172, n174, n175, n178, n181, n182, n186, n188,
         n190, n192, n193, n194, n195, n198, n199, n201, n202, n204, n205,
         n206, n207, n208, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U6 ( .A(n3), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U8 ( .A(n4), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U10 ( .A(n370), .B(n5), .Z(DIFF[9]) );
  XOR2_X1 U42 ( .A(n74), .B(n334), .Z(DIFF[48]) );
  XOR2_X1 U43 ( .A(n335), .B(n352), .Z(DIFF[49]) );
  XOR2_X1 U44 ( .A(n15), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U45 ( .A(n9), .B(n336), .Z(DIFF[50]) );
  XOR2_X1 U46 ( .A(n12), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U47 ( .A(n16), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U49 ( .A(n64), .B(n338), .Z(DIFF[52]) );
  XOR2_X1 U50 ( .A(n339), .B(n353), .Z(DIFF[53]) );
  XOR2_X1 U51 ( .A(n10), .B(n340), .Z(DIFF[54]) );
  XOR2_X1 U59 ( .A(n43), .B(B[61]), .Z(DIFF[61]) );
  XOR2_X1 U60 ( .A(n40), .B(n347), .Z(DIFF[62]) );
  XOR2_X1 U61 ( .A(n343), .B(n354), .Z(DIFF[57]) );
  XOR2_X1 U71 ( .A(n55), .B(n342), .Z(DIFF[56]) );
  XOR2_X1 U72 ( .A(n11), .B(n344), .Z(DIFF[58]) );
  XOR2_X1 U73 ( .A(n45), .B(n346), .Z(DIFF[60]) );
  XOR2_X1 U90 ( .A(n160), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U96 ( .A(n350), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U100 ( .A(n92), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U101 ( .A(n112), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n311), .B(n151), .Z(DIFF[25]) );
  XOR2_X1 U113 ( .A(n306), .B(n349), .Z(DIFF[20]) );
  XOR2_X1 U123 ( .A(n312), .B(n150), .Z(DIFF[26]) );
  XOR2_X1 U127 ( .A(n316), .B(n139), .Z(DIFF[30]) );
  XOR2_X1 U128 ( .A(n314), .B(n143), .Z(DIFF[28]) );
  XOR2_X1 U129 ( .A(n310), .B(n14), .Z(DIFF[24]) );
  XOR2_X1 U130 ( .A(n162), .B(n302), .Z(DIFF[16]) );
  XOR2_X1 U131 ( .A(n315), .B(n140), .Z(DIFF[29]) );
  XOR2_X1 U132 ( .A(n123), .B(n320), .Z(DIFF[34]) );
  XOR2_X1 U133 ( .A(n303), .B(n20), .Z(DIFF[17]) );
  XOR2_X1 U134 ( .A(n308), .B(n159), .Z(DIFF[22]) );
  XOR2_X1 U135 ( .A(n304), .B(n21), .Z(DIFF[18]) );
  XOR2_X1 U146 ( .A(n111), .B(n324), .Z(DIFF[38]) );
  XOR2_X1 U153 ( .A(n322), .B(n351), .Z(DIFF[36]) );
  XOR2_X1 U154 ( .A(n319), .B(n124), .Z(DIFF[33]) );
  XOR2_X1 U199 ( .A(n362), .B(n28), .Z(DIFF[2]) );
  XOR2_X1 U200 ( .A(n364), .B(n359), .Z(DIFF[4]) );
  XOR2_X1 U201 ( .A(n368), .B(n8), .Z(DIFF[8]) );
  XOR2_X1 U202 ( .A(n366), .B(n39), .Z(DIFF[5]) );
  XOR2_X1 U204 ( .A(n367), .B(n36), .Z(DIFF[6]) );
  NAND3_X1 U227 ( .A1(n344), .A2(n345), .A3(n343), .ZN(n48) );
  NAND3_X1 U228 ( .A1(n340), .A2(n341), .A3(n339), .ZN(n58) );
  NAND3_X1 U229 ( .A1(n336), .A2(n337), .A3(n335), .ZN(n67) );
  NAND3_X1 U230 ( .A1(n357), .A2(n22), .A3(n79), .ZN(n77) );
  NAND3_X1 U245 ( .A1(n356), .A2(n19), .A3(n130), .ZN(n128) );
  NAND3_X1 U250 ( .A1(n359), .A2(n297), .A3(n178), .ZN(n175) );
  NAND3_X1 U254 ( .A1(n181), .A2(n27), .A3(n182), .ZN(n174) );
  NAND3_X1 U258 ( .A1(n299), .A2(n300), .A3(n1), .ZN(n186) );
  NAND3_X1 U267 ( .A1(n369), .A2(n359), .A3(n27), .ZN(n199) );
  XOR2_X1 U5 ( .A(n300), .B(n204), .Z(DIFF[14]) );
  XOR2_X1 U9 ( .A(B[7]), .B(n205), .Z(DIFF[7]) );
  XOR2_X1 U55 ( .A(n206), .B(B[63]), .Z(DIFF[63]) );
  INV_X1 U3 ( .A(n57), .ZN(n353) );
  INV_X1 U4 ( .A(n47), .ZN(n354) );
  NOR2_X1 U7 ( .A1(n12), .A2(B[45]), .ZN(n88) );
  XNOR2_X1 U11 ( .A(n337), .B(n71), .ZN(DIFF[51]) );
  NAND2_X1 U12 ( .A1(n336), .A2(n9), .ZN(n71) );
  AND2_X1 U13 ( .A1(n335), .A2(n352), .ZN(n9) );
  INV_X1 U14 ( .A(n66), .ZN(n352) );
  NOR2_X1 U15 ( .A1(n66), .A2(n67), .ZN(n64) );
  NOR2_X1 U16 ( .A1(n57), .A2(n58), .ZN(n55) );
  NOR2_X1 U17 ( .A1(n47), .A2(n48), .ZN(n45) );
  XNOR2_X1 U18 ( .A(n341), .B(n62), .ZN(DIFF[55]) );
  NAND2_X1 U19 ( .A1(n340), .A2(n10), .ZN(n62) );
  XNOR2_X1 U20 ( .A(n345), .B(n53), .ZN(DIFF[59]) );
  NAND2_X1 U21 ( .A1(n344), .A2(n11), .ZN(n53) );
  NAND2_X1 U22 ( .A1(n64), .A2(n338), .ZN(n57) );
  NAND2_X1 U23 ( .A1(n55), .A2(n342), .ZN(n47) );
  NAND2_X1 U24 ( .A1(n45), .A2(n346), .ZN(n43) );
  AND2_X1 U25 ( .A1(n339), .A2(n353), .ZN(n10) );
  AND2_X1 U26 ( .A1(n343), .A2(n354), .ZN(n11) );
  NAND2_X1 U27 ( .A1(n330), .A2(n331), .ZN(n81) );
  INV_X1 U28 ( .A(n14), .ZN(n348) );
  NAND2_X1 U29 ( .A1(n328), .A2(n98), .ZN(n3) );
  NOR2_X1 U30 ( .A1(n15), .A2(B[41]), .ZN(n98) );
  XNOR2_X1 U31 ( .A(n98), .B(B[42]), .ZN(DIFF[42]) );
  XNOR2_X1 U32 ( .A(n88), .B(B[46]), .ZN(DIFF[46]) );
  NAND2_X1 U33 ( .A1(n74), .A2(n334), .ZN(n66) );
  OR2_X1 U34 ( .A1(n16), .A2(B[44]), .ZN(n12) );
  INV_X1 U35 ( .A(n114), .ZN(n350) );
  NAND2_X1 U36 ( .A1(n332), .A2(n88), .ZN(n4) );
  NAND2_X1 U37 ( .A1(n40), .A2(n347), .ZN(n206) );
  NOR2_X1 U38 ( .A1(B[61]), .A2(n43), .ZN(n40) );
  NAND2_X1 U39 ( .A1(n332), .A2(n333), .ZN(n80) );
  NOR2_X1 U40 ( .A1(n160), .A2(B[21]), .ZN(n159) );
  NOR2_X1 U41 ( .A1(n348), .A2(n137), .ZN(n143) );
  XNOR2_X1 U48 ( .A(n138), .B(n317), .ZN(DIFF[31]) );
  NAND2_X1 U52 ( .A1(n139), .A2(n316), .ZN(n138) );
  INV_X1 U53 ( .A(n127), .ZN(n349) );
  AND2_X1 U54 ( .A1(n19), .A2(n349), .ZN(n14) );
  AND2_X1 U56 ( .A1(n140), .A2(n315), .ZN(n139) );
  NOR2_X1 U57 ( .A1(n127), .A2(n128), .ZN(n114) );
  NOR2_X1 U58 ( .A1(n131), .A2(n132), .ZN(n130) );
  INV_X1 U62 ( .A(n137), .ZN(n356) );
  NOR2_X1 U63 ( .A1(n112), .A2(B[37]), .ZN(n111) );
  NOR2_X1 U64 ( .A1(n76), .A2(n77), .ZN(n74) );
  NOR2_X1 U65 ( .A1(n80), .A2(n81), .ZN(n79) );
  INV_X1 U66 ( .A(n86), .ZN(n357) );
  NOR2_X1 U67 ( .A1(B[32]), .A2(n350), .ZN(n124) );
  INV_X1 U68 ( .A(n76), .ZN(n351) );
  NAND2_X1 U69 ( .A1(n22), .A2(n351), .ZN(n92) );
  OR2_X1 U70 ( .A1(B[40]), .A2(n92), .ZN(n15) );
  NAND2_X1 U74 ( .A1(n316), .A2(n317), .ZN(n131) );
  OR2_X1 U75 ( .A1(n92), .A2(n86), .ZN(n16) );
  NOR2_X1 U76 ( .A1(n188), .A2(n360), .ZN(n204) );
  NAND2_X1 U77 ( .A1(n355), .A2(n190), .ZN(n188) );
  NOR2_X1 U78 ( .A1(B[12]), .A2(n298), .ZN(n190) );
  XNOR2_X1 U79 ( .A(n301), .B(n186), .ZN(DIFF[15]) );
  XNOR2_X1 U80 ( .A(n1), .B(n298), .ZN(DIFF[13]) );
  NAND2_X1 U81 ( .A1(n349), .A2(n306), .ZN(n160) );
  NAND2_X1 U82 ( .A1(n162), .A2(n163), .ZN(n127) );
  NOR2_X1 U83 ( .A1(n164), .A2(n165), .ZN(n163) );
  NAND2_X1 U84 ( .A1(n302), .A2(n305), .ZN(n164) );
  NAND2_X1 U85 ( .A1(n303), .A2(n304), .ZN(n165) );
  INV_X1 U86 ( .A(B[12]), .ZN(n297) );
  INV_X1 U87 ( .A(n194), .ZN(n355) );
  XNOR2_X1 U88 ( .A(n313), .B(n149), .ZN(DIFF[27]) );
  NAND2_X1 U89 ( .A1(n312), .A2(n150), .ZN(n149) );
  XNOR2_X1 U91 ( .A(n309), .B(n158), .ZN(DIFF[23]) );
  NAND2_X1 U92 ( .A1(n308), .A2(n159), .ZN(n158) );
  AND2_X1 U93 ( .A1(n151), .A2(n311), .ZN(n150) );
  AND3_X1 U94 ( .A1(n302), .A2(n301), .A3(n172), .ZN(n20) );
  AND2_X1 U95 ( .A1(n301), .A2(n172), .ZN(n162) );
  AND2_X1 U97 ( .A1(n303), .A2(n20), .ZN(n21) );
  AND2_X1 U98 ( .A1(n143), .A2(n314), .ZN(n140) );
  AND4_X1 U99 ( .A1(n306), .A2(n309), .A3(n308), .A4(n307), .ZN(n19) );
  XNOR2_X1 U102 ( .A(n294), .B(n305), .ZN(DIFF[19]) );
  NAND2_X1 U103 ( .A1(n21), .A2(n304), .ZN(n294) );
  NAND4_X1 U104 ( .A1(n310), .A2(n313), .A3(n312), .A4(n311), .ZN(n137) );
  NAND4_X1 U105 ( .A1(n326), .A2(n329), .A3(n328), .A4(n327), .ZN(n86) );
  XNOR2_X1 U107 ( .A(n208), .B(n321), .ZN(DIFF[35]) );
  NAND2_X1 U108 ( .A1(n320), .A2(n123), .ZN(n208) );
  NAND2_X1 U109 ( .A1(n114), .A2(n115), .ZN(n76) );
  NOR2_X1 U110 ( .A1(n116), .A2(n117), .ZN(n115) );
  NAND2_X1 U111 ( .A1(n319), .A2(n320), .ZN(n117) );
  NAND2_X1 U112 ( .A1(n318), .A2(n321), .ZN(n116) );
  NAND2_X1 U114 ( .A1(n351), .A2(n322), .ZN(n112) );
  AND2_X1 U115 ( .A1(n124), .A2(n319), .ZN(n123) );
  XNOR2_X1 U116 ( .A(n207), .B(n325), .ZN(DIFF[39]) );
  NAND2_X1 U117 ( .A1(n324), .A2(n111), .ZN(n207) );
  NAND2_X1 U118 ( .A1(n314), .A2(n315), .ZN(n132) );
  AND4_X1 U119 ( .A1(n322), .A2(n325), .A3(n324), .A4(n323), .ZN(n22) );
  NAND4_X1 U120 ( .A1(n370), .A2(n368), .A3(n296), .A4(n295), .ZN(n194) );
  NOR2_X1 U121 ( .A1(B[24]), .A2(n348), .ZN(n151) );
  XNOR2_X1 U122 ( .A(n24), .B(B[11]), .ZN(DIFF[11]) );
  NOR2_X1 U124 ( .A1(n25), .A2(n26), .ZN(n24) );
  OR2_X1 U125 ( .A1(n365), .A2(n198), .ZN(n26) );
  OR2_X1 U126 ( .A1(B[10]), .A2(n73), .ZN(n25) );
  NOR2_X1 U136 ( .A1(n174), .A2(n175), .ZN(n172) );
  NOR2_X1 U137 ( .A1(B[10]), .A2(B[11]), .ZN(n178) );
  NOR2_X1 U138 ( .A1(B[14]), .A2(n298), .ZN(n182) );
  AND2_X1 U139 ( .A1(n192), .A2(n8), .ZN(n1) );
  NOR2_X1 U140 ( .A1(n194), .A2(B[12]), .ZN(n192) );
  INV_X1 U141 ( .A(n73), .ZN(n359) );
  XNOR2_X1 U142 ( .A(n363), .B(n107), .ZN(DIFF[3]) );
  NAND2_X1 U143 ( .A1(n362), .A2(n28), .ZN(n107) );
  AND2_X1 U144 ( .A1(n39), .A2(n366), .ZN(n36) );
  INV_X1 U145 ( .A(n8), .ZN(n360) );
  AND2_X1 U147 ( .A1(n364), .A2(n359), .ZN(n39) );
  INV_X1 U148 ( .A(n27), .ZN(n365) );
  XNOR2_X1 U149 ( .A(n297), .B(n195), .ZN(DIFF[12]) );
  NAND2_X1 U150 ( .A1(n2), .A2(n355), .ZN(n195) );
  AND3_X1 U151 ( .A1(n359), .A2(n363), .A3(n27), .ZN(n2) );
  XNOR2_X1 U152 ( .A(n199), .B(n295), .ZN(DIFF[10]) );
  INV_X1 U155 ( .A(n198), .ZN(n369) );
  NOR2_X1 U156 ( .A1(n360), .A2(B[8]), .ZN(n5) );
  NAND2_X1 U157 ( .A1(n367), .A2(n36), .ZN(n205) );
  AND2_X1 U158 ( .A1(n6), .A2(n7), .ZN(n27) );
  NOR2_X1 U159 ( .A1(B[5]), .A2(B[4]), .ZN(n6) );
  NOR2_X1 U160 ( .A1(B[7]), .A2(B[6]), .ZN(n7) );
  NAND2_X1 U161 ( .A1(n201), .A2(n202), .ZN(n73) );
  NOR2_X1 U162 ( .A1(B[1]), .A2(\B[0] ), .ZN(n201) );
  NOR2_X1 U163 ( .A1(B[3]), .A2(B[2]), .ZN(n202) );
  AND2_X1 U164 ( .A1(n193), .A2(n27), .ZN(n8) );
  NOR2_X1 U165 ( .A1(n73), .A2(B[3]), .ZN(n193) );
  INV_X1 U166 ( .A(B[1]), .ZN(n361) );
  AND2_X1 U167 ( .A1(n361), .A2(n358), .ZN(n28) );
  INV_X1 U168 ( .A(\B[0] ), .ZN(n358) );
  INV_X1 U169 ( .A(B[3]), .ZN(n363) );
  INV_X1 U170 ( .A(B[8]), .ZN(n368) );
  INV_X1 U171 ( .A(B[6]), .ZN(n367) );
  INV_X1 U172 ( .A(B[2]), .ZN(n362) );
  INV_X1 U173 ( .A(B[9]), .ZN(n370) );
  OR2_X1 U174 ( .A1(B[9]), .A2(B[8]), .ZN(n198) );
  INV_X1 U175 ( .A(B[5]), .ZN(n366) );
  INV_X1 U176 ( .A(B[4]), .ZN(n364) );
  XNOR2_X1 U177 ( .A(\B[0] ), .B(n361), .ZN(DIFF[1]) );
  NOR2_X1 U178 ( .A1(B[9]), .A2(B[8]), .ZN(n181) );
  INV_X1 U179 ( .A(B[10]), .ZN(n295) );
  INV_X1 U180 ( .A(B[11]), .ZN(n296) );
  INV_X1 U181 ( .A(n299), .ZN(n298) );
  INV_X1 U182 ( .A(B[13]), .ZN(n299) );
  INV_X1 U183 ( .A(B[14]), .ZN(n300) );
  INV_X1 U184 ( .A(B[15]), .ZN(n301) );
  INV_X1 U185 ( .A(B[16]), .ZN(n302) );
  INV_X1 U186 ( .A(B[17]), .ZN(n303) );
  INV_X1 U187 ( .A(B[18]), .ZN(n304) );
  INV_X1 U188 ( .A(B[19]), .ZN(n305) );
  INV_X1 U189 ( .A(B[20]), .ZN(n306) );
  INV_X1 U190 ( .A(B[21]), .ZN(n307) );
  INV_X1 U191 ( .A(B[22]), .ZN(n308) );
  INV_X1 U192 ( .A(B[23]), .ZN(n309) );
  INV_X1 U193 ( .A(B[24]), .ZN(n310) );
  INV_X1 U194 ( .A(B[25]), .ZN(n311) );
  INV_X1 U195 ( .A(B[26]), .ZN(n312) );
  INV_X1 U196 ( .A(B[27]), .ZN(n313) );
  INV_X1 U197 ( .A(B[28]), .ZN(n314) );
  INV_X1 U198 ( .A(B[29]), .ZN(n315) );
  INV_X1 U203 ( .A(B[30]), .ZN(n316) );
  INV_X1 U205 ( .A(B[31]), .ZN(n317) );
  INV_X1 U206 ( .A(B[32]), .ZN(n318) );
  INV_X1 U207 ( .A(B[33]), .ZN(n319) );
  INV_X1 U208 ( .A(B[34]), .ZN(n320) );
  INV_X1 U209 ( .A(B[35]), .ZN(n321) );
  INV_X1 U210 ( .A(B[36]), .ZN(n322) );
  INV_X1 U211 ( .A(B[37]), .ZN(n323) );
  INV_X1 U212 ( .A(B[38]), .ZN(n324) );
  INV_X1 U213 ( .A(B[39]), .ZN(n325) );
  INV_X1 U214 ( .A(B[40]), .ZN(n326) );
  INV_X1 U215 ( .A(B[41]), .ZN(n327) );
  INV_X1 U216 ( .A(B[42]), .ZN(n328) );
  INV_X1 U217 ( .A(B[43]), .ZN(n329) );
  INV_X1 U218 ( .A(B[44]), .ZN(n330) );
  INV_X1 U219 ( .A(B[45]), .ZN(n331) );
  INV_X1 U220 ( .A(B[46]), .ZN(n332) );
  INV_X1 U221 ( .A(B[47]), .ZN(n333) );
  INV_X1 U222 ( .A(B[48]), .ZN(n334) );
  INV_X1 U223 ( .A(B[49]), .ZN(n335) );
  INV_X1 U224 ( .A(B[50]), .ZN(n336) );
  INV_X1 U225 ( .A(B[51]), .ZN(n337) );
  INV_X1 U226 ( .A(B[52]), .ZN(n338) );
  INV_X1 U231 ( .A(B[53]), .ZN(n339) );
  INV_X1 U232 ( .A(B[54]), .ZN(n340) );
  INV_X1 U233 ( .A(B[55]), .ZN(n341) );
  INV_X1 U234 ( .A(B[56]), .ZN(n342) );
  INV_X1 U235 ( .A(B[57]), .ZN(n343) );
  INV_X1 U236 ( .A(B[58]), .ZN(n344) );
  INV_X1 U237 ( .A(B[59]), .ZN(n345) );
  INV_X1 U238 ( .A(B[60]), .ZN(n346) );
  INV_X1 U239 ( .A(B[62]), .ZN(n347) );
endmodule


module complement_NBIT64_22 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_22_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_21_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n228, n229, n230, n231, n232, n234, n235, n237, n238, n239,
         n240, n242, n243, n244, n246, n247, n248, n250, n251, n252, n254,
         n255, n256, n257, n258, n260, n261, n262, n264, n265, n266, n267,
         n268, n270, n271, n272, n274, n275, n276, n278, n279, n280, n281,
         n282, n284, n285, n286, n287, n288, n289, n290, n291, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U113 ( .A(n228), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U114 ( .A(n230), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U116 ( .A(n234), .B(B[62]), .Z(DIFF[62]) );
  NAND3_X1 U117 ( .A1(n315), .A2(n316), .A3(n235), .ZN(n234) );
  XOR2_X1 U119 ( .A(n237), .B(B[58]), .Z(DIFF[58]) );
  NAND3_X1 U120 ( .A1(n313), .A2(n314), .A3(n240), .ZN(n237) );
  XOR2_X1 U122 ( .A(n242), .B(B[54]), .Z(DIFF[54]) );
  NAND3_X1 U123 ( .A1(n311), .A2(n312), .A3(n244), .ZN(n242) );
  XOR2_X1 U125 ( .A(n246), .B(B[50]), .Z(DIFF[50]) );
  NAND3_X1 U126 ( .A1(n309), .A2(n310), .A3(n248), .ZN(n246) );
  XOR2_X1 U127 ( .A(n232), .B(B[4]), .Z(DIFF[4]) );
  XOR2_X1 U129 ( .A(n250), .B(B[46]), .Z(DIFF[46]) );
  NAND3_X1 U130 ( .A1(n307), .A2(n308), .A3(n252), .ZN(n250) );
  XOR2_X1 U132 ( .A(n254), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U133 ( .A(n256), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U135 ( .A(n261), .B(B[38]), .Z(DIFF[38]) );
  NAND3_X1 U136 ( .A1(n303), .A2(n304), .A3(n262), .ZN(n261) );
  XOR2_X1 U138 ( .A(n264), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U139 ( .A(n266), .B(B[32]), .Z(DIFF[32]) );
  NAND3_X1 U140 ( .A1(n300), .A2(n301), .A3(n268), .ZN(n266) );
  XOR2_X1 U142 ( .A(n260), .B(B[2]), .Z(DIFF[2]) );
  XOR2_X1 U143 ( .A(n270), .B(B[28]), .Z(DIFF[28]) );
  NAND3_X1 U144 ( .A1(n298), .A2(n299), .A3(n272), .ZN(n270) );
  XOR2_X1 U146 ( .A(n274), .B(B[24]), .Z(DIFF[24]) );
  NAND3_X1 U147 ( .A1(n296), .A2(n297), .A3(n276), .ZN(n274) );
  XOR2_X1 U149 ( .A(n278), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U150 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U151 ( .A(n281), .B(B[18]), .Z(DIFF[18]) );
  NAND3_X1 U152 ( .A1(n293), .A2(n294), .A3(n282), .ZN(n281) );
  XOR2_X1 U154 ( .A(n284), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U155 ( .A(n287), .B(B[12]), .Z(DIFF[12]) );
  NAND3_X1 U156 ( .A1(n229), .A2(n319), .A3(n288), .ZN(n287) );
  XOR2_X1 U157 ( .A(n289), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U43 ( .A(n295), .B(n280), .Z(DIFF[19]) );
  XOR2_X1 U52 ( .A(n302), .B(n265), .Z(DIFF[34]) );
  XOR2_X1 U54 ( .A(n210), .B(n304), .Z(DIFF[37]) );
  XOR2_X1 U56 ( .A(n292), .B(n286), .Z(DIFF[13]) );
  XOR2_X1 U57 ( .A(n306), .B(n255), .Z(DIFF[42]) );
  XOR2_X1 U58 ( .A(n305), .B(n258), .Z(DIFF[39]) );
  NOR3_X1 U3 ( .A1(B[50]), .A2(B[51]), .A3(n246), .ZN(n244) );
  NOR3_X1 U4 ( .A1(B[54]), .A2(B[55]), .A3(n242), .ZN(n240) );
  NOR3_X1 U5 ( .A1(B[58]), .A2(B[59]), .A3(n237), .ZN(n235) );
  NOR3_X1 U6 ( .A1(B[46]), .A2(B[47]), .A3(n250), .ZN(n248) );
  NOR2_X1 U7 ( .A1(n254), .A2(B[43]), .ZN(n252) );
  NOR2_X1 U8 ( .A1(n264), .A2(B[35]), .ZN(n262) );
  NAND2_X1 U9 ( .A1(n280), .A2(n295), .ZN(n278) );
  NAND2_X1 U10 ( .A1(n286), .A2(n292), .ZN(n284) );
  NAND2_X1 U11 ( .A1(n258), .A2(n305), .ZN(n256) );
  NAND2_X1 U12 ( .A1(n265), .A2(n302), .ZN(n264) );
  NAND2_X1 U13 ( .A1(n255), .A2(n306), .ZN(n254) );
  NOR3_X1 U14 ( .A1(B[14]), .A2(B[15]), .A3(n284), .ZN(n282) );
  NOR3_X1 U15 ( .A1(B[24]), .A2(B[25]), .A3(n274), .ZN(n272) );
  NOR3_X1 U16 ( .A1(B[28]), .A2(B[29]), .A3(n270), .ZN(n268) );
  NOR3_X1 U17 ( .A1(B[20]), .A2(B[21]), .A3(n278), .ZN(n276) );
  NOR3_X1 U18 ( .A1(B[32]), .A2(B[33]), .A3(n266), .ZN(n265) );
  NOR3_X1 U19 ( .A1(B[40]), .A2(B[41]), .A3(n256), .ZN(n255) );
  NAND2_X1 U20 ( .A1(n290), .A2(n319), .ZN(n289) );
  NOR2_X1 U21 ( .A1(n281), .A2(B[18]), .ZN(n280) );
  NOR2_X1 U22 ( .A1(n261), .A2(B[38]), .ZN(n258) );
  XNOR2_X1 U23 ( .A(B[16]), .B(n282), .ZN(DIFF[16]) );
  XNOR2_X1 U24 ( .A(n206), .B(n294), .ZN(DIFF[17]) );
  NAND2_X1 U25 ( .A1(n282), .A2(n293), .ZN(n206) );
  XNOR2_X1 U26 ( .A(n208), .B(n297), .ZN(DIFF[23]) );
  NAND2_X1 U27 ( .A1(n276), .A2(n296), .ZN(n208) );
  XNOR2_X1 U28 ( .A(B[21]), .B(n279), .ZN(DIFF[21]) );
  NOR2_X1 U29 ( .A1(B[20]), .A2(n278), .ZN(n279) );
  XNOR2_X1 U30 ( .A(B[22]), .B(n276), .ZN(DIFF[22]) );
  XNOR2_X1 U31 ( .A(n207), .B(n299), .ZN(DIFF[27]) );
  NAND2_X1 U32 ( .A1(n272), .A2(n298), .ZN(n207) );
  XNOR2_X1 U33 ( .A(n205), .B(n301), .ZN(DIFF[31]) );
  NAND2_X1 U34 ( .A1(n268), .A2(n300), .ZN(n205) );
  XNOR2_X1 U35 ( .A(B[29]), .B(n271), .ZN(DIFF[29]) );
  NOR2_X1 U36 ( .A1(B[28]), .A2(n270), .ZN(n271) );
  XNOR2_X1 U37 ( .A(B[30]), .B(n268), .ZN(DIFF[30]) );
  XNOR2_X1 U38 ( .A(B[41]), .B(n257), .ZN(DIFF[41]) );
  NOR2_X1 U39 ( .A1(B[40]), .A2(n256), .ZN(n257) );
  AND2_X1 U40 ( .A1(n262), .A2(n303), .ZN(n210) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n262), .ZN(DIFF[36]) );
  XNOR2_X1 U42 ( .A(n201), .B(n308), .ZN(DIFF[45]) );
  NAND2_X1 U44 ( .A1(n252), .A2(n307), .ZN(n201) );
  XNOR2_X1 U45 ( .A(B[47]), .B(n251), .ZN(DIFF[47]) );
  NOR2_X1 U46 ( .A1(B[46]), .A2(n250), .ZN(n251) );
  XNOR2_X1 U47 ( .A(B[44]), .B(n252), .ZN(DIFF[44]) );
  XNOR2_X1 U48 ( .A(B[48]), .B(n248), .ZN(DIFF[48]) );
  XNOR2_X1 U49 ( .A(n200), .B(n310), .ZN(DIFF[49]) );
  NAND2_X1 U50 ( .A1(n248), .A2(n309), .ZN(n200) );
  XNOR2_X1 U51 ( .A(B[51]), .B(n247), .ZN(DIFF[51]) );
  NOR2_X1 U53 ( .A1(B[50]), .A2(n246), .ZN(n247) );
  XNOR2_X1 U55 ( .A(B[52]), .B(n244), .ZN(DIFF[52]) );
  XNOR2_X1 U59 ( .A(n202), .B(n312), .ZN(DIFF[53]) );
  NAND2_X1 U60 ( .A1(n244), .A2(n311), .ZN(n202) );
  XNOR2_X1 U61 ( .A(B[56]), .B(n240), .ZN(DIFF[56]) );
  XNOR2_X1 U62 ( .A(n203), .B(n314), .ZN(DIFF[57]) );
  NAND2_X1 U63 ( .A1(n240), .A2(n313), .ZN(n203) );
  XNOR2_X1 U64 ( .A(n204), .B(n316), .ZN(DIFF[61]) );
  NAND2_X1 U65 ( .A1(n235), .A2(n315), .ZN(n204) );
  XNOR2_X1 U66 ( .A(n209), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U67 ( .A1(n234), .A2(B[62]), .ZN(n209) );
  XNOR2_X1 U68 ( .A(B[59]), .B(n239), .ZN(DIFF[59]) );
  NOR2_X1 U69 ( .A1(B[58]), .A2(n237), .ZN(n239) );
  XNOR2_X1 U70 ( .A(B[60]), .B(n235), .ZN(DIFF[60]) );
  XNOR2_X1 U71 ( .A(B[15]), .B(n285), .ZN(DIFF[15]) );
  NOR2_X1 U72 ( .A1(B[14]), .A2(n284), .ZN(n285) );
  XNOR2_X1 U73 ( .A(B[25]), .B(n275), .ZN(DIFF[25]) );
  NOR2_X1 U74 ( .A1(B[24]), .A2(n274), .ZN(n275) );
  XNOR2_X1 U75 ( .A(B[33]), .B(n267), .ZN(DIFF[33]) );
  NOR2_X1 U76 ( .A1(B[32]), .A2(n266), .ZN(n267) );
  XNOR2_X1 U77 ( .A(B[55]), .B(n243), .ZN(DIFF[55]) );
  NOR2_X1 U78 ( .A1(B[54]), .A2(n242), .ZN(n243) );
  XNOR2_X1 U79 ( .A(B[26]), .B(n272), .ZN(DIFF[26]) );
  NOR3_X1 U80 ( .A1(B[11]), .A2(B[9]), .A3(B[8]), .ZN(n288) );
  NOR3_X1 U81 ( .A1(n232), .A2(B[4]), .A3(n291), .ZN(n229) );
  OR3_X1 U82 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n291) );
  NOR3_X1 U83 ( .A1(B[4]), .A2(B[5]), .A3(n232), .ZN(n231) );
  NOR2_X1 U84 ( .A1(n228), .A2(B[9]), .ZN(n290) );
  XNOR2_X1 U85 ( .A(B[6]), .B(n231), .ZN(DIFF[6]) );
  XNOR2_X1 U86 ( .A(n229), .B(B[8]), .ZN(DIFF[8]) );
  NAND2_X1 U87 ( .A1(n231), .A2(n317), .ZN(n230) );
  INV_X1 U88 ( .A(B[6]), .ZN(n317) );
  XNOR2_X1 U89 ( .A(B[5]), .B(n238), .ZN(DIFF[5]) );
  NOR2_X1 U90 ( .A1(B[4]), .A2(n232), .ZN(n238) );
  XNOR2_X1 U91 ( .A(n211), .B(B[3]), .ZN(DIFF[3]) );
  NOR2_X1 U92 ( .A1(n260), .A2(B[2]), .ZN(n211) );
  XNOR2_X1 U93 ( .A(n290), .B(B[10]), .ZN(DIFF[10]) );
  NAND2_X1 U94 ( .A1(n229), .A2(n318), .ZN(n228) );
  INV_X1 U95 ( .A(B[8]), .ZN(n318) );
  OR3_X1 U96 ( .A1(B[2]), .A2(B[3]), .A3(n260), .ZN(n232) );
  OR2_X1 U97 ( .A1(B[1]), .A2(\B[0] ), .ZN(n260) );
  INV_X1 U98 ( .A(B[10]), .ZN(n319) );
  NOR2_X1 U99 ( .A1(n287), .A2(B[12]), .ZN(n286) );
  INV_X1 U100 ( .A(B[13]), .ZN(n292) );
  INV_X1 U101 ( .A(B[16]), .ZN(n293) );
  INV_X1 U102 ( .A(B[17]), .ZN(n294) );
  INV_X1 U103 ( .A(B[19]), .ZN(n295) );
  INV_X1 U104 ( .A(B[22]), .ZN(n296) );
  INV_X1 U105 ( .A(B[23]), .ZN(n297) );
  INV_X1 U106 ( .A(B[26]), .ZN(n298) );
  INV_X1 U107 ( .A(B[27]), .ZN(n299) );
  INV_X1 U108 ( .A(B[30]), .ZN(n300) );
  INV_X1 U109 ( .A(B[31]), .ZN(n301) );
  INV_X1 U110 ( .A(B[34]), .ZN(n302) );
  INV_X1 U111 ( .A(B[36]), .ZN(n303) );
  INV_X1 U112 ( .A(B[37]), .ZN(n304) );
  INV_X1 U115 ( .A(B[39]), .ZN(n305) );
  INV_X1 U118 ( .A(B[42]), .ZN(n306) );
  INV_X1 U121 ( .A(B[44]), .ZN(n307) );
  INV_X1 U124 ( .A(B[45]), .ZN(n308) );
  INV_X1 U128 ( .A(B[48]), .ZN(n309) );
  INV_X1 U131 ( .A(B[49]), .ZN(n310) );
  INV_X1 U134 ( .A(B[52]), .ZN(n311) );
  INV_X1 U137 ( .A(B[53]), .ZN(n312) );
  INV_X1 U141 ( .A(B[56]), .ZN(n313) );
  INV_X1 U145 ( .A(B[57]), .ZN(n314) );
  INV_X1 U148 ( .A(B[60]), .ZN(n315) );
  INV_X1 U153 ( .A(B[61]), .ZN(n316) );
endmodule


module complement_NBIT64_21 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_21_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_20_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n19, n20, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n86, n90, n93, n95, n96, n98,
         n99, n100, n105, n106, n107, n108, n110, n114, n115, n116, n117, n119,
         n123, n125, n126, n127, n128, n129, n130, n131, n132, n135, n137,
         n138, n141, n142, n143, n144, n150, n152, n153, n156, n157, n158,
         n159, n160, n161, n162, n163, n168, n170, n171, n174, n175, n176,
         n177, n180, n182, n183, n188, n189, n190, n192, n193, n196, n197,
         n198, n199, n201, n203, n204, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U13 ( .A(n326), .B(n4), .Z(DIFF[51]) );
  XOR2_X1 U20 ( .A(n323), .B(n5), .Z(DIFF[47]) );
  XOR2_X1 U22 ( .A(n329), .B(n6), .Z(DIFF[55]) );
  XOR2_X1 U27 ( .A(n303), .B(n7), .Z(DIFF[15]) );
  XOR2_X1 U31 ( .A(n308), .B(n8), .Z(DIFF[23]) );
  XOR2_X1 U33 ( .A(n301), .B(n9), .Z(DIFF[12]) );
  XOR2_X1 U35 ( .A(n310), .B(n10), .Z(DIFF[27]) );
  XOR2_X1 U37 ( .A(n313), .B(n11), .Z(DIFF[31]) );
  XOR2_X1 U41 ( .A(n306), .B(n12), .Z(DIFF[19]) );
  XOR2_X1 U43 ( .A(n320), .B(n13), .Z(DIFF[43]) );
  XOR2_X1 U45 ( .A(n318), .B(n14), .Z(DIFF[39]) );
  XOR2_X1 U47 ( .A(n316), .B(n15), .Z(DIFF[35]) );
  XOR2_X1 U3 ( .A(B[59]), .B(n212), .Z(DIFF[59]) );
  XOR2_X1 U5 ( .A(n302), .B(n213), .Z(DIFF[13]) );
  XOR2_X1 U7 ( .A(B[3]), .B(n214), .Z(DIFF[3]) );
  XOR2_X1 U54 ( .A(n114), .B(n327), .Z(DIFF[52]) );
  XOR2_X1 U58 ( .A(n105), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U61 ( .A(n332), .B(n95), .Z(DIFF[61]) );
  XOR2_X1 U62 ( .A(n96), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U76 ( .A(n324), .B(n28), .Z(DIFF[48]) );
  XOR2_X1 U137 ( .A(B[20]), .B(n163), .Z(DIFF[20]) );
  XOR2_X1 U150 ( .A(B[36]), .B(n132), .Z(DIFF[36]) );
  XOR2_X1 U194 ( .A(n123), .B(B[4]), .Z(DIFF[4]) );
  XNOR2_X1 U4 ( .A(B[58]), .B(n19), .ZN(DIFF[58]) );
  INV_X1 U6 ( .A(n108), .ZN(n341) );
  AND2_X1 U8 ( .A1(n339), .A2(n325), .ZN(n119) );
  AND2_X1 U9 ( .A1(n330), .A2(n342), .ZN(n19) );
  AND2_X1 U10 ( .A1(n95), .A2(n332), .ZN(n93) );
  AND2_X1 U11 ( .A1(n341), .A2(n328), .ZN(n110) );
  NAND2_X1 U12 ( .A1(n327), .A2(n114), .ZN(n108) );
  INV_X1 U14 ( .A(n100), .ZN(n342) );
  XNOR2_X1 U15 ( .A(B[46]), .B(n20), .ZN(DIFF[46]) );
  XNOR2_X1 U16 ( .A(B[50]), .B(n119), .ZN(DIFF[50]) );
  XNOR2_X1 U17 ( .A(B[45]), .B(n23), .ZN(DIFF[45]) );
  XNOR2_X1 U18 ( .A(B[49]), .B(n339), .ZN(DIFF[49]) );
  XNOR2_X1 U19 ( .A(B[33]), .B(n34), .ZN(DIFF[33]) );
  NOR2_X1 U21 ( .A1(n345), .A2(B[46]), .ZN(n5) );
  INV_X1 U23 ( .A(n20), .ZN(n345) );
  NOR2_X1 U24 ( .A1(n338), .A2(B[50]), .ZN(n4) );
  INV_X1 U25 ( .A(n119), .ZN(n338) );
  AND2_X1 U26 ( .A1(n322), .A2(n23), .ZN(n20) );
  INV_X1 U28 ( .A(n116), .ZN(n339) );
  NOR2_X1 U29 ( .A1(n115), .A2(n116), .ZN(n114) );
  NAND2_X1 U30 ( .A1(n117), .A2(n325), .ZN(n115) );
  NOR2_X1 U32 ( .A1(B[51]), .A2(B[50]), .ZN(n117) );
  XNOR2_X1 U34 ( .A(B[54]), .B(n110), .ZN(DIFF[54]) );
  XNOR2_X1 U36 ( .A(B[53]), .B(n341), .ZN(DIFF[53]) );
  XNOR2_X1 U38 ( .A(B[57]), .B(n342), .ZN(DIFF[57]) );
  XNOR2_X1 U39 ( .A(B[62]), .B(n93), .ZN(DIFF[62]) );
  NOR2_X1 U40 ( .A1(n96), .A2(B[60]), .ZN(n95) );
  XNOR2_X1 U42 ( .A(B[63]), .B(n217), .ZN(DIFF[63]) );
  NOR2_X1 U44 ( .A1(n343), .A2(B[62]), .ZN(n217) );
  INV_X1 U46 ( .A(n93), .ZN(n343) );
  NOR2_X1 U48 ( .A1(n340), .A2(B[54]), .ZN(n6) );
  INV_X1 U49 ( .A(n110), .ZN(n340) );
  OR2_X1 U50 ( .A1(n100), .A2(n98), .ZN(n96) );
  NAND2_X1 U51 ( .A1(n99), .A2(n330), .ZN(n98) );
  NOR2_X1 U52 ( .A1(B[59]), .A2(B[58]), .ZN(n99) );
  NAND2_X1 U53 ( .A1(n131), .A2(n322), .ZN(n130) );
  NOR2_X1 U55 ( .A1(B[47]), .A2(B[46]), .ZN(n131) );
  OR2_X1 U56 ( .A1(B[56]), .A2(n105), .ZN(n100) );
  OR2_X1 U57 ( .A1(n108), .A2(n106), .ZN(n105) );
  NAND2_X1 U59 ( .A1(n107), .A2(n328), .ZN(n106) );
  NOR2_X1 U60 ( .A1(B[55]), .A2(B[54]), .ZN(n107) );
  NAND2_X1 U63 ( .A1(n331), .A2(n19), .ZN(n212) );
  NOR2_X1 U64 ( .A1(n352), .A2(n192), .ZN(n7) );
  NAND2_X1 U65 ( .A1(n193), .A2(n27), .ZN(n192) );
  NOR2_X1 U66 ( .A1(B[14]), .A2(B[13]), .ZN(n193) );
  AND2_X1 U67 ( .A1(n305), .A2(n26), .ZN(n24) );
  AND2_X1 U68 ( .A1(n304), .A2(n1), .ZN(n26) );
  INV_X1 U69 ( .A(n175), .ZN(n336) );
  NOR2_X1 U70 ( .A1(n352), .A2(n349), .ZN(n213) );
  INV_X1 U71 ( .A(n27), .ZN(n349) );
  XNOR2_X1 U72 ( .A(B[37]), .B(n150), .ZN(DIFF[37]) );
  XNOR2_X1 U73 ( .A(B[32]), .B(n29), .ZN(DIFF[32]) );
  XNOR2_X1 U74 ( .A(B[28]), .B(n168), .ZN(DIFF[28]) );
  XNOR2_X1 U75 ( .A(B[44]), .B(n135), .ZN(DIFF[44]) );
  AND2_X1 U77 ( .A1(n312), .A2(n31), .ZN(n25) );
  AND2_X1 U78 ( .A1(n315), .A2(n34), .ZN(n37) );
  NAND2_X1 U79 ( .A1(n324), .A2(n28), .ZN(n116) );
  AND2_X1 U80 ( .A1(n314), .A2(n29), .ZN(n34) );
  AND2_X1 U81 ( .A1(n321), .A2(n135), .ZN(n23) );
  INV_X1 U82 ( .A(n142), .ZN(n346) );
  INV_X1 U83 ( .A(n30), .ZN(n352) );
  NOR2_X1 U84 ( .A1(n163), .A2(n160), .ZN(n175) );
  XNOR2_X1 U85 ( .A(B[25]), .B(n174), .ZN(DIFF[25]) );
  XNOR2_X1 U86 ( .A(B[21]), .B(n180), .ZN(DIFF[21]) );
  AND2_X1 U87 ( .A1(n309), .A2(n174), .ZN(n33) );
  AND2_X1 U88 ( .A1(n307), .A2(n180), .ZN(n32) );
  AND4_X1 U89 ( .A1(n357), .A2(n359), .A3(n353), .A4(n188), .ZN(n1) );
  AND2_X1 U90 ( .A1(n189), .A2(n190), .ZN(n188) );
  NOR2_X1 U91 ( .A1(B[13]), .A2(n300), .ZN(n189) );
  NOR2_X1 U92 ( .A1(B[15]), .A2(B[14]), .ZN(n190) );
  AND2_X1 U93 ( .A1(n359), .A2(n301), .ZN(n27) );
  NAND2_X1 U94 ( .A1(n197), .A2(n359), .ZN(n16) );
  NOR2_X1 U95 ( .A1(B[13]), .A2(n300), .ZN(n197) );
  NOR2_X1 U96 ( .A1(n163), .A2(n156), .ZN(n29) );
  NAND2_X1 U97 ( .A1(n157), .A2(n158), .ZN(n156) );
  NOR2_X1 U98 ( .A1(n160), .A2(n161), .ZN(n157) );
  NOR2_X1 U99 ( .A1(B[28]), .A2(n159), .ZN(n158) );
  NOR2_X1 U100 ( .A1(n132), .A2(n129), .ZN(n142) );
  NOR2_X1 U101 ( .A1(n132), .A2(B[36]), .ZN(n150) );
  NOR2_X1 U102 ( .A1(n336), .A2(n159), .ZN(n168) );
  NOR2_X1 U103 ( .A1(n346), .A2(n128), .ZN(n135) );
  NOR2_X1 U104 ( .A1(n132), .A2(n125), .ZN(n28) );
  NAND2_X1 U105 ( .A1(n126), .A2(n127), .ZN(n125) );
  NOR2_X1 U106 ( .A1(n129), .A2(n130), .ZN(n126) );
  NOR2_X1 U107 ( .A1(B[44]), .A2(n128), .ZN(n127) );
  XNOR2_X1 U108 ( .A(B[29]), .B(n31), .ZN(DIFF[29]) );
  XNOR2_X1 U109 ( .A(B[41]), .B(n141), .ZN(DIFF[41]) );
  AND2_X1 U110 ( .A1(n319), .A2(n141), .ZN(n36) );
  AND2_X1 U111 ( .A1(n317), .A2(n150), .ZN(n35) );
  AND2_X1 U112 ( .A1(n311), .A2(n168), .ZN(n31) );
  AND2_X1 U113 ( .A1(n357), .A2(n353), .ZN(n30) );
  NOR2_X1 U114 ( .A1(n348), .A2(B[22]), .ZN(n8) );
  INV_X1 U115 ( .A(n32), .ZN(n348) );
  NOR2_X1 U116 ( .A1(n336), .A2(B[24]), .ZN(n174) );
  NOR2_X1 U117 ( .A1(n163), .A2(B[20]), .ZN(n180) );
  NAND2_X1 U118 ( .A1(n2), .A2(n1), .ZN(n163) );
  AND2_X1 U119 ( .A1(n182), .A2(n183), .ZN(n2) );
  NOR2_X1 U120 ( .A1(B[19]), .A2(B[18]), .ZN(n183) );
  NOR2_X1 U121 ( .A1(B[17]), .A2(B[16]), .ZN(n182) );
  XNOR2_X1 U122 ( .A(B[26]), .B(n33), .ZN(DIFF[26]) );
  XNOR2_X1 U123 ( .A(B[22]), .B(n32), .ZN(DIFF[22]) );
  NOR2_X1 U124 ( .A1(n334), .A2(B[26]), .ZN(n10) );
  INV_X1 U125 ( .A(n33), .ZN(n334) );
  NOR2_X1 U126 ( .A1(n337), .A2(B[34]), .ZN(n15) );
  INV_X1 U127 ( .A(n37), .ZN(n337) );
  NOR2_X1 U128 ( .A1(n346), .A2(B[40]), .ZN(n141) );
  NAND2_X1 U129 ( .A1(n3), .A2(n29), .ZN(n132) );
  AND2_X1 U130 ( .A1(n152), .A2(n153), .ZN(n3) );
  NOR2_X1 U131 ( .A1(B[35]), .A2(B[34]), .ZN(n153) );
  NOR2_X1 U132 ( .A1(B[33]), .A2(B[32]), .ZN(n152) );
  XNOR2_X1 U133 ( .A(B[42]), .B(n36), .ZN(DIFF[42]) );
  XNOR2_X1 U134 ( .A(B[40]), .B(n142), .ZN(DIFF[40]) );
  XNOR2_X1 U135 ( .A(B[24]), .B(n175), .ZN(DIFF[24]) );
  XNOR2_X1 U136 ( .A(B[38]), .B(n35), .ZN(DIFF[38]) );
  XNOR2_X1 U138 ( .A(B[30]), .B(n25), .ZN(DIFF[30]) );
  XNOR2_X1 U139 ( .A(B[34]), .B(n37), .ZN(DIFF[34]) );
  NOR2_X1 U140 ( .A1(n344), .A2(B[42]), .ZN(n13) );
  INV_X1 U141 ( .A(n36), .ZN(n344) );
  NOR2_X1 U142 ( .A1(n347), .A2(B[38]), .ZN(n14) );
  INV_X1 U143 ( .A(n35), .ZN(n347) );
  NOR2_X1 U144 ( .A1(n335), .A2(B[30]), .ZN(n11) );
  INV_X1 U145 ( .A(n25), .ZN(n335) );
  NAND2_X1 U146 ( .A1(n170), .A2(n171), .ZN(n159) );
  NOR2_X1 U147 ( .A1(B[27]), .A2(B[26]), .ZN(n171) );
  NOR2_X1 U148 ( .A1(B[25]), .A2(B[24]), .ZN(n170) );
  NAND2_X1 U149 ( .A1(n176), .A2(n177), .ZN(n160) );
  NOR2_X1 U151 ( .A1(B[23]), .A2(B[22]), .ZN(n177) );
  NOR2_X1 U152 ( .A1(B[21]), .A2(B[20]), .ZN(n176) );
  NAND2_X1 U153 ( .A1(n143), .A2(n144), .ZN(n129) );
  NOR2_X1 U154 ( .A1(B[39]), .A2(B[38]), .ZN(n144) );
  NOR2_X1 U155 ( .A1(B[37]), .A2(B[36]), .ZN(n143) );
  NAND2_X1 U156 ( .A1(n162), .A2(n312), .ZN(n161) );
  NOR2_X1 U157 ( .A1(B[31]), .A2(B[30]), .ZN(n162) );
  NAND2_X1 U158 ( .A1(n137), .A2(n138), .ZN(n128) );
  NOR2_X1 U159 ( .A1(B[41]), .A2(B[40]), .ZN(n137) );
  NOR2_X1 U160 ( .A1(B[43]), .A2(B[42]), .ZN(n138) );
  INV_X1 U161 ( .A(n201), .ZN(n359) );
  INV_X1 U162 ( .A(n123), .ZN(n353) );
  INV_X1 U163 ( .A(n199), .ZN(n357) );
  NOR2_X1 U164 ( .A1(n352), .A2(n201), .ZN(n9) );
  XNOR2_X1 U165 ( .A(B[17]), .B(n26), .ZN(DIFF[17]) );
  XNOR2_X1 U166 ( .A(B[18]), .B(n24), .ZN(DIFF[18]) );
  XNOR2_X1 U167 ( .A(B[16]), .B(n1), .ZN(DIFF[16]) );
  XNOR2_X1 U168 ( .A(n196), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U169 ( .A1(n198), .A2(n16), .ZN(n196) );
  OR2_X1 U170 ( .A1(n199), .A2(n123), .ZN(n198) );
  NOR2_X1 U171 ( .A1(n333), .A2(B[18]), .ZN(n12) );
  INV_X1 U172 ( .A(n24), .ZN(n333) );
  NAND2_X1 U173 ( .A1(n356), .A2(n38), .ZN(n214) );
  INV_X1 U174 ( .A(B[2]), .ZN(n356) );
  NOR2_X1 U175 ( .A1(n352), .A2(B[8]), .ZN(n86) );
  NOR2_X1 U176 ( .A1(n123), .A2(B[4]), .ZN(n90) );
  NAND2_X1 U177 ( .A1(n208), .A2(n209), .ZN(n123) );
  NOR2_X1 U178 ( .A1(B[1]), .A2(\B[0] ), .ZN(n208) );
  NOR2_X1 U179 ( .A1(B[3]), .A2(B[2]), .ZN(n209) );
  XNOR2_X1 U180 ( .A(B[5]), .B(n90), .ZN(DIFF[5]) );
  XNOR2_X1 U181 ( .A(B[9]), .B(n86), .ZN(DIFF[9]) );
  XNOR2_X1 U182 ( .A(B[8]), .B(n30), .ZN(DIFF[8]) );
  XNOR2_X1 U183 ( .A(B[6]), .B(n39), .ZN(DIFF[6]) );
  XNOR2_X1 U184 ( .A(B[10]), .B(n40), .ZN(DIFF[10]) );
  XNOR2_X1 U185 ( .A(B[2]), .B(n38), .ZN(DIFF[2]) );
  XNOR2_X1 U186 ( .A(B[7]), .B(n215), .ZN(DIFF[7]) );
  NOR2_X1 U187 ( .A1(n354), .A2(B[6]), .ZN(n215) );
  INV_X1 U188 ( .A(n39), .ZN(n354) );
  XNOR2_X1 U189 ( .A(B[11]), .B(n216), .ZN(DIFF[11]) );
  NOR2_X1 U190 ( .A1(n351), .A2(B[10]), .ZN(n216) );
  INV_X1 U191 ( .A(n40), .ZN(n351) );
  AND2_X1 U192 ( .A1(n358), .A2(n90), .ZN(n39) );
  INV_X1 U193 ( .A(B[5]), .ZN(n358) );
  AND2_X1 U195 ( .A1(n360), .A2(n86), .ZN(n40) );
  INV_X1 U196 ( .A(B[9]), .ZN(n360) );
  NAND2_X1 U197 ( .A1(n203), .A2(n204), .ZN(n201) );
  NOR2_X1 U198 ( .A1(B[11]), .A2(B[10]), .ZN(n203) );
  NOR2_X1 U199 ( .A1(B[9]), .A2(B[8]), .ZN(n204) );
  NAND2_X1 U200 ( .A1(n210), .A2(n211), .ZN(n199) );
  NOR2_X1 U201 ( .A1(B[5]), .A2(B[4]), .ZN(n210) );
  NOR2_X1 U202 ( .A1(B[7]), .A2(B[6]), .ZN(n211) );
  AND2_X1 U203 ( .A1(n355), .A2(n350), .ZN(n38) );
  INV_X1 U204 ( .A(\B[0] ), .ZN(n350) );
  INV_X1 U205 ( .A(B[1]), .ZN(n355) );
  XNOR2_X1 U206 ( .A(n355), .B(\B[0] ), .ZN(DIFF[1]) );
  INV_X1 U207 ( .A(n301), .ZN(n300) );
  INV_X1 U208 ( .A(B[12]), .ZN(n301) );
  INV_X1 U209 ( .A(B[13]), .ZN(n302) );
  INV_X1 U210 ( .A(B[15]), .ZN(n303) );
  INV_X1 U211 ( .A(B[16]), .ZN(n304) );
  INV_X1 U212 ( .A(B[17]), .ZN(n305) );
  INV_X1 U213 ( .A(B[19]), .ZN(n306) );
  INV_X1 U214 ( .A(B[21]), .ZN(n307) );
  INV_X1 U215 ( .A(B[23]), .ZN(n308) );
  INV_X1 U216 ( .A(B[25]), .ZN(n309) );
  INV_X1 U217 ( .A(B[27]), .ZN(n310) );
  INV_X1 U218 ( .A(B[28]), .ZN(n311) );
  INV_X1 U219 ( .A(B[29]), .ZN(n312) );
  INV_X1 U220 ( .A(B[31]), .ZN(n313) );
  INV_X1 U221 ( .A(B[32]), .ZN(n314) );
  INV_X1 U222 ( .A(B[33]), .ZN(n315) );
  INV_X1 U223 ( .A(B[35]), .ZN(n316) );
  INV_X1 U224 ( .A(B[37]), .ZN(n317) );
  INV_X1 U225 ( .A(B[39]), .ZN(n318) );
  INV_X1 U226 ( .A(B[41]), .ZN(n319) );
  INV_X1 U227 ( .A(B[43]), .ZN(n320) );
  INV_X1 U228 ( .A(B[44]), .ZN(n321) );
  INV_X1 U229 ( .A(B[45]), .ZN(n322) );
  INV_X1 U230 ( .A(B[47]), .ZN(n323) );
  INV_X1 U231 ( .A(B[48]), .ZN(n324) );
  INV_X1 U232 ( .A(B[49]), .ZN(n325) );
  INV_X1 U233 ( .A(B[51]), .ZN(n326) );
  INV_X1 U234 ( .A(B[52]), .ZN(n327) );
  INV_X1 U235 ( .A(B[53]), .ZN(n328) );
  INV_X1 U236 ( .A(B[55]), .ZN(n329) );
  INV_X1 U237 ( .A(B[57]), .ZN(n330) );
  INV_X1 U238 ( .A(B[58]), .ZN(n331) );
  INV_X1 U239 ( .A(B[61]), .ZN(n332) );
endmodule


module complement_NBIT64_20 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_20_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_19_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n210, n211, n212, n214, n215, n216, n218, n219, n220, n222,
         n223, n224, n226, n227, n228, n229, n231, n232, n233, n234, n235,
         n237, n238, n239, n240, n242, n243, n244, n246, n247, n248, n249,
         n250, n251, n252, n254, n255, n256, n257, n258, n259, n260, n261,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U96 ( .A(n199), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U97 ( .A(n201), .B(B[6]), .Z(DIFF[6]) );
  NAND3_X1 U98 ( .A1(n268), .A2(n269), .A3(n202), .ZN(n201) );
  XOR2_X1 U99 ( .A(n203), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U100 ( .A(n205), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U101 ( .A(n208), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U103 ( .A(n207), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U104 ( .A(n210), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U106 ( .A(n212), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U107 ( .A(n214), .B(B[52]), .Z(DIFF[52]) );
  XOR2_X1 U109 ( .A(n216), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U110 ( .A(n218), .B(B[48]), .Z(DIFF[48]) );
  XOR2_X1 U112 ( .A(n220), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U113 ( .A(n222), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U115 ( .A(n224), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U116 ( .A(n226), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U117 ( .A(n229), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U119 ( .A(n228), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U120 ( .A(n231), .B(B[36]), .Z(DIFF[36]) );
  XOR2_X1 U121 ( .A(n234), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U123 ( .A(n235), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U124 ( .A(n237), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U126 ( .A(n239), .B(B[28]), .Z(DIFF[28]) );
  XOR2_X1 U127 ( .A(n242), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U129 ( .A(n244), .B(B[24]), .Z(DIFF[24]) );
  XOR2_X1 U130 ( .A(n246), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U131 ( .A(n248), .B(B[20]), .Z(DIFF[20]) );
  XOR2_X1 U132 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U133 ( .A(n251), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U135 ( .A(n252), .B(B[16]), .Z(DIFF[16]) );
  XOR2_X1 U136 ( .A(n254), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U137 ( .A(n256), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U138 ( .A(n260), .B(B[10]), .Z(DIFF[10]) );
  NAND3_X1 U139 ( .A1(n202), .A2(n268), .A3(n261), .ZN(n199) );
  XOR2_X1 U20 ( .A(n204), .B(n266), .Z(DIFF[62]) );
  XOR2_X1 U27 ( .A(n265), .B(n233), .Z(DIFF[35]) );
  XOR2_X1 U33 ( .A(n255), .B(n262), .Z(DIFF[14]) );
  XOR2_X1 U35 ( .A(n247), .B(n264), .Z(DIFF[22]) );
  XOR2_X1 U39 ( .A(n263), .B(n250), .Z(DIFF[19]) );
  NOR3_X1 U3 ( .A1(B[60]), .A2(B[61]), .A3(n205), .ZN(n204) );
  OR3_X1 U4 ( .A1(B[58]), .A2(B[59]), .A3(n207), .ZN(n205) );
  OR3_X1 U5 ( .A1(B[50]), .A2(B[51]), .A3(n216), .ZN(n214) );
  OR3_X1 U6 ( .A1(B[54]), .A2(B[55]), .A3(n212), .ZN(n210) );
  OR3_X1 U7 ( .A1(B[48]), .A2(B[49]), .A3(n218), .ZN(n216) );
  OR3_X1 U8 ( .A1(B[52]), .A2(B[53]), .A3(n214), .ZN(n212) );
  OR3_X1 U9 ( .A1(B[56]), .A2(B[57]), .A3(n210), .ZN(n207) );
  OR3_X1 U10 ( .A1(B[46]), .A2(B[47]), .A3(n220), .ZN(n218) );
  NOR2_X1 U11 ( .A1(n251), .A2(B[18]), .ZN(n250) );
  NOR2_X1 U12 ( .A1(n234), .A2(B[34]), .ZN(n233) );
  NAND2_X1 U13 ( .A1(n233), .A2(n265), .ZN(n231) );
  NAND2_X1 U14 ( .A1(n250), .A2(n263), .ZN(n248) );
  OR2_X1 U15 ( .A1(n254), .A2(B[15]), .ZN(n252) );
  OR3_X1 U16 ( .A1(B[32]), .A2(B[33]), .A3(n235), .ZN(n234) );
  NAND2_X1 U17 ( .A1(n247), .A2(n264), .ZN(n246) );
  OR3_X1 U18 ( .A1(B[44]), .A2(B[45]), .A3(n222), .ZN(n220) );
  NAND2_X1 U19 ( .A1(n255), .A2(n262), .ZN(n254) );
  NOR3_X1 U21 ( .A1(B[20]), .A2(B[21]), .A3(n248), .ZN(n247) );
  XNOR2_X1 U22 ( .A(n194), .B(B[17]), .ZN(DIFF[17]) );
  NOR2_X1 U23 ( .A1(n252), .A2(B[16]), .ZN(n194) );
  NOR2_X1 U24 ( .A1(n256), .A2(B[13]), .ZN(n255) );
  OR2_X1 U25 ( .A1(n246), .A2(B[23]), .ZN(n244) );
  OR3_X1 U26 ( .A1(B[28]), .A2(B[29]), .A3(n239), .ZN(n237) );
  OR3_X1 U28 ( .A1(B[42]), .A2(B[43]), .A3(n224), .ZN(n222) );
  OR3_X1 U29 ( .A1(B[24]), .A2(B[25]), .A3(n244), .ZN(n242) );
  OR3_X1 U30 ( .A1(B[38]), .A2(B[39]), .A3(n228), .ZN(n226) );
  OR3_X1 U31 ( .A1(B[30]), .A2(B[31]), .A3(n237), .ZN(n235) );
  OR3_X1 U32 ( .A1(B[40]), .A2(B[41]), .A3(n226), .ZN(n224) );
  OR3_X1 U34 ( .A1(B[26]), .A2(B[27]), .A3(n242), .ZN(n239) );
  OR3_X1 U36 ( .A1(B[36]), .A2(B[37]), .A3(n231), .ZN(n228) );
  OR3_X1 U37 ( .A1(B[16]), .A2(B[17]), .A3(n252), .ZN(n251) );
  NAND2_X1 U38 ( .A1(n204), .A2(n266), .ZN(n203) );
  XNOR2_X1 U40 ( .A(n197), .B(B[25]), .ZN(DIFF[25]) );
  NOR2_X1 U41 ( .A1(n244), .A2(B[24]), .ZN(n197) );
  XNOR2_X1 U42 ( .A(B[21]), .B(n249), .ZN(DIFF[21]) );
  NOR2_X1 U43 ( .A1(B[20]), .A2(n248), .ZN(n249) );
  XNOR2_X1 U44 ( .A(B[27]), .B(n243), .ZN(DIFF[27]) );
  NOR2_X1 U45 ( .A1(B[26]), .A2(n242), .ZN(n243) );
  XNOR2_X1 U46 ( .A(B[31]), .B(n238), .ZN(DIFF[31]) );
  NOR2_X1 U47 ( .A1(B[30]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U48 ( .A(n193), .B(B[29]), .ZN(DIFF[29]) );
  NOR2_X1 U49 ( .A1(n239), .A2(B[28]), .ZN(n193) );
  XNOR2_X1 U50 ( .A(n192), .B(B[33]), .ZN(DIFF[33]) );
  NOR2_X1 U51 ( .A1(n235), .A2(B[32]), .ZN(n192) );
  XNOR2_X1 U52 ( .A(B[37]), .B(n232), .ZN(DIFF[37]) );
  NOR2_X1 U53 ( .A1(B[36]), .A2(n231), .ZN(n232) );
  XNOR2_X1 U54 ( .A(n195), .B(B[39]), .ZN(DIFF[39]) );
  NOR2_X1 U55 ( .A1(n228), .A2(B[38]), .ZN(n195) );
  XNOR2_X1 U56 ( .A(B[41]), .B(n227), .ZN(DIFF[41]) );
  NOR2_X1 U57 ( .A1(B[40]), .A2(n226), .ZN(n227) );
  XNOR2_X1 U58 ( .A(n196), .B(B[43]), .ZN(DIFF[43]) );
  NOR2_X1 U59 ( .A1(n224), .A2(B[42]), .ZN(n196) );
  XNOR2_X1 U60 ( .A(B[45]), .B(n223), .ZN(DIFF[45]) );
  NOR2_X1 U61 ( .A1(B[44]), .A2(n222), .ZN(n223) );
  XNOR2_X1 U62 ( .A(n191), .B(B[47]), .ZN(DIFF[47]) );
  NOR2_X1 U63 ( .A1(n220), .A2(B[46]), .ZN(n191) );
  XNOR2_X1 U64 ( .A(n188), .B(B[51]), .ZN(DIFF[51]) );
  NOR2_X1 U65 ( .A1(n216), .A2(B[50]), .ZN(n188) );
  XNOR2_X1 U66 ( .A(B[49]), .B(n219), .ZN(DIFF[49]) );
  NOR2_X1 U67 ( .A1(B[48]), .A2(n218), .ZN(n219) );
  XNOR2_X1 U68 ( .A(B[53]), .B(n215), .ZN(DIFF[53]) );
  NOR2_X1 U69 ( .A1(B[52]), .A2(n214), .ZN(n215) );
  XNOR2_X1 U70 ( .A(n189), .B(B[55]), .ZN(DIFF[55]) );
  NOR2_X1 U71 ( .A1(n212), .A2(B[54]), .ZN(n189) );
  XNOR2_X1 U72 ( .A(B[57]), .B(n211), .ZN(DIFF[57]) );
  NOR2_X1 U73 ( .A1(B[56]), .A2(n210), .ZN(n211) );
  XNOR2_X1 U74 ( .A(n190), .B(B[59]), .ZN(DIFF[59]) );
  NOR2_X1 U75 ( .A1(n207), .A2(B[58]), .ZN(n190) );
  XNOR2_X1 U76 ( .A(B[61]), .B(n206), .ZN(DIFF[61]) );
  NOR2_X1 U77 ( .A1(B[60]), .A2(n205), .ZN(n206) );
  NOR3_X1 U78 ( .A1(n199), .A2(B[10]), .A3(n258), .ZN(n257) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[9]), .A3(B[8]), .ZN(n258) );
  NOR2_X1 U80 ( .A1(n229), .A2(B[3]), .ZN(n202) );
  NOR3_X1 U81 ( .A1(B[5]), .A2(B[7]), .A3(B[6]), .ZN(n261) );
  NOR2_X1 U82 ( .A1(n199), .A2(B[8]), .ZN(n198) );
  INV_X1 U83 ( .A(B[5]), .ZN(n269) );
  XNOR2_X1 U84 ( .A(n202), .B(B[4]), .ZN(DIFF[4]) );
  NAND2_X1 U85 ( .A1(n202), .A2(n268), .ZN(n208) );
  XNOR2_X1 U86 ( .A(B[9]), .B(n198), .ZN(DIFF[9]) );
  XNOR2_X1 U87 ( .A(B[7]), .B(n200), .ZN(DIFF[7]) );
  NOR2_X1 U88 ( .A1(B[6]), .A2(n201), .ZN(n200) );
  XNOR2_X1 U89 ( .A(B[11]), .B(n259), .ZN(DIFF[11]) );
  NOR2_X1 U90 ( .A1(B[10]), .A2(n260), .ZN(n259) );
  XNOR2_X1 U91 ( .A(n240), .B(B[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U92 ( .A(n257), .B(B[12]), .ZN(DIFF[12]) );
  NAND2_X1 U93 ( .A1(n257), .A2(n271), .ZN(n256) );
  INV_X1 U94 ( .A(B[12]), .ZN(n271) );
  NAND2_X1 U95 ( .A1(n198), .A2(n270), .ZN(n260) );
  INV_X1 U102 ( .A(B[9]), .ZN(n270) );
  NAND2_X1 U105 ( .A1(n240), .A2(n267), .ZN(n229) );
  INV_X1 U108 ( .A(B[2]), .ZN(n267) );
  INV_X1 U111 ( .A(B[4]), .ZN(n268) );
  NOR2_X1 U114 ( .A1(B[1]), .A2(\B[0] ), .ZN(n240) );
  INV_X1 U118 ( .A(B[14]), .ZN(n262) );
  INV_X1 U122 ( .A(B[19]), .ZN(n263) );
  INV_X1 U125 ( .A(B[22]), .ZN(n264) );
  INV_X1 U128 ( .A(B[35]), .ZN(n265) );
  INV_X1 U134 ( .A(B[62]), .ZN(n266) );
endmodule


module complement_NBIT64_19 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_19_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_18_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32,
         n34, n38, n41, n44, n46, n48, n49, n54, n56, n58, n59, n63, n65, n67,
         n68, n72, n74, n76, n77, n80, n81, n82, n87, n88, n89, n90, n92, n97,
         n98, n110, n112, n114, n115, n116, n121, n122, n123, n126, n130, n131,
         n132, n133, n134, n139, n140, n141, n144, n150, n151, n152, n153,
         n158, n159, n167, n172, n177, n178, n179, n181, n182, n183, n184,
         n187, n188, n189, n192, n193, n195, n196, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U8 ( .A(n5), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U10 ( .A(n6), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U15 ( .A(n289), .B(n9), .Z(DIFF[14]) );
  XOR2_X1 U17 ( .A(n361), .B(n10), .Z(DIFF[12]) );
  XOR2_X1 U27 ( .A(n16), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U45 ( .A(n322), .B(n90), .Z(DIFF[46]) );
  XOR2_X1 U48 ( .A(n74), .B(n324), .Z(DIFF[48]) );
  XOR2_X1 U49 ( .A(n19), .B(n334), .Z(DIFF[58]) );
  XOR2_X1 U50 ( .A(n325), .B(n342), .Z(DIFF[49]) );
  XOR2_X1 U51 ( .A(n329), .B(n343), .Z(DIFF[53]) );
  XOR2_X1 U52 ( .A(n333), .B(n344), .Z(DIFF[57]) );
  XOR2_X1 U59 ( .A(n17), .B(n326), .Z(DIFF[50]) );
  XOR2_X1 U60 ( .A(n65), .B(n328), .Z(DIFF[52]) );
  XOR2_X1 U61 ( .A(n18), .B(n330), .Z(DIFF[54]) );
  XOR2_X1 U65 ( .A(n56), .B(n332), .Z(DIFF[56]) );
  XOR2_X1 U66 ( .A(n46), .B(n336), .Z(DIFF[60]) );
  XOR2_X1 U78 ( .A(n41), .B(n337), .Z(DIFF[62]) );
  XOR2_X1 U79 ( .A(n44), .B(B[61]), .Z(DIFF[61]) );
  XOR2_X1 U91 ( .A(n22), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U94 ( .A(n112), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U97 ( .A(n21), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U98 ( .A(n1), .B(n320), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n340), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U118 ( .A(n301), .B(n151), .Z(DIFF[26]) );
  XOR2_X1 U133 ( .A(n305), .B(n140), .Z(DIFF[30]) );
  XOR2_X1 U134 ( .A(n304), .B(n141), .Z(DIFF[29]) );
  XOR2_X1 U135 ( .A(n303), .B(n144), .Z(DIFF[28]) );
  XOR2_X1 U139 ( .A(n296), .B(n2), .Z(DIFF[21]) );
  XOR2_X1 U140 ( .A(n300), .B(n26), .Z(DIFF[25]) );
  XOR2_X1 U141 ( .A(n122), .B(n309), .Z(DIFF[34]) );
  XOR2_X1 U142 ( .A(n297), .B(n159), .Z(DIFF[22]) );
  XOR2_X1 U143 ( .A(n299), .B(n23), .Z(DIFF[24]) );
  XOR2_X1 U144 ( .A(n308), .B(n123), .Z(DIFF[33]) );
  XOR2_X1 U145 ( .A(n311), .B(n341), .Z(DIFF[36]) );
  XOR2_X1 U146 ( .A(n317), .B(n98), .Z(DIFF[42]) );
  XOR2_X1 U147 ( .A(n319), .B(n92), .Z(DIFF[44]) );
  XOR2_X1 U206 ( .A(n357), .B(n29), .Z(DIFF[5]) );
  XOR2_X1 U207 ( .A(n355), .B(n352), .Z(DIFF[4]) );
  XOR2_X1 U208 ( .A(n28), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U211 ( .A(n358), .B(n38), .Z(DIFF[6]) );
  XOR2_X1 U213 ( .A(n360), .B(n199), .Z(DIFF[10]) );
  NAND3_X1 U238 ( .A1(n334), .A2(n335), .A3(n333), .ZN(n49) );
  NAND3_X1 U239 ( .A1(n330), .A2(n331), .A3(n329), .ZN(n59) );
  NAND3_X1 U240 ( .A1(n326), .A2(n327), .A3(n325), .ZN(n68) );
  NAND3_X1 U241 ( .A1(n349), .A2(n348), .A3(n80), .ZN(n77) );
  NAND3_X1 U262 ( .A1(n362), .A2(n361), .A3(n31), .ZN(n192) );
  XOR2_X1 U3 ( .A(n202), .B(B[15]), .Z(DIFF[15]) );
  NAND3_X1 U4 ( .A1(n187), .A2(n352), .A3(n188), .ZN(n202) );
  XOR2_X1 U9 ( .A(B[7]), .B(n205), .Z(DIFF[7]) );
  XOR2_X1 U46 ( .A(n207), .B(B[63]), .Z(DIFF[63]) );
  INV_X1 U5 ( .A(n58), .ZN(n343) );
  INV_X1 U6 ( .A(n48), .ZN(n344) );
  NOR2_X1 U7 ( .A1(n67), .A2(n68), .ZN(n65) );
  NOR2_X1 U11 ( .A1(n58), .A2(n59), .ZN(n56) );
  NOR2_X1 U12 ( .A1(n48), .A2(n49), .ZN(n46) );
  NAND2_X1 U13 ( .A1(n65), .A2(n328), .ZN(n58) );
  NAND2_X1 U14 ( .A1(n56), .A2(n332), .ZN(n48) );
  NAND2_X1 U16 ( .A1(n46), .A2(n336), .ZN(n44) );
  AND2_X1 U18 ( .A1(n325), .A2(n342), .ZN(n17) );
  AND2_X1 U19 ( .A1(n329), .A2(n343), .ZN(n18) );
  AND2_X1 U20 ( .A1(n333), .A2(n344), .ZN(n19) );
  INV_X1 U21 ( .A(n67), .ZN(n342) );
  INV_X1 U22 ( .A(n4), .ZN(n340) );
  NOR2_X1 U23 ( .A1(B[61]), .A2(n44), .ZN(n41) );
  NAND2_X1 U24 ( .A1(n74), .A2(n324), .ZN(n67) );
  NOR2_X1 U25 ( .A1(n112), .A2(B[37]), .ZN(n110) );
  NAND4_X1 U26 ( .A1(n290), .A2(n294), .A3(n293), .A4(n292), .ZN(n153) );
  NOR2_X1 U28 ( .A1(n1), .A2(n320), .ZN(n90) );
  NOR2_X1 U29 ( .A1(n22), .A2(B[41]), .ZN(n98) );
  NOR2_X1 U30 ( .A1(n21), .A2(n88), .ZN(n92) );
  NOR2_X1 U31 ( .A1(n339), .A2(n131), .ZN(n144) );
  INV_X1 U32 ( .A(n23), .ZN(n339) );
  NOR2_X1 U33 ( .A1(B[32]), .A2(n340), .ZN(n123) );
  INV_X1 U34 ( .A(B[14]), .ZN(n289) );
  OR2_X1 U35 ( .A1(n76), .A2(n87), .ZN(n21) );
  AND2_X1 U36 ( .A1(n26), .A2(n300), .ZN(n151) );
  AND2_X1 U37 ( .A1(n123), .A2(n308), .ZN(n122) );
  AND4_X1 U38 ( .A1(n126), .A2(n346), .A3(n347), .A4(n345), .ZN(n4) );
  INV_X1 U39 ( .A(n131), .ZN(n347) );
  NOR2_X1 U40 ( .A1(n133), .A2(n134), .ZN(n126) );
  INV_X1 U41 ( .A(n132), .ZN(n346) );
  AND2_X1 U42 ( .A1(n141), .A2(n304), .ZN(n140) );
  OR2_X1 U43 ( .A1(B[40]), .A2(n21), .ZN(n22) );
  INV_X1 U44 ( .A(n76), .ZN(n341) );
  INV_X1 U47 ( .A(n130), .ZN(n345) );
  NOR2_X1 U53 ( .A1(n76), .A2(n77), .ZN(n74) );
  INV_X1 U54 ( .A(n88), .ZN(n349) );
  INV_X1 U55 ( .A(n87), .ZN(n348) );
  NAND2_X1 U56 ( .A1(n167), .A2(n209), .ZN(n5) );
  NOR3_X1 U57 ( .A1(B[16]), .A2(n291), .A3(B[18]), .ZN(n167) );
  NAND2_X1 U58 ( .A1(n172), .A2(n209), .ZN(n6) );
  NOR2_X1 U62 ( .A1(n291), .A2(B[16]), .ZN(n172) );
  NOR2_X1 U63 ( .A1(n24), .A2(n152), .ZN(n23) );
  OR2_X1 U64 ( .A1(n132), .A2(n153), .ZN(n24) );
  NOR3_X1 U67 ( .A1(B[15]), .A2(n288), .A3(n356), .ZN(n8) );
  NAND4_X1 U68 ( .A1(n299), .A2(n302), .A3(n301), .A4(n300), .ZN(n131) );
  NAND4_X1 U69 ( .A1(n295), .A2(n298), .A3(n297), .A4(n296), .ZN(n132) );
  NAND2_X1 U70 ( .A1(n4), .A2(n114), .ZN(n76) );
  NOR2_X1 U71 ( .A1(n115), .A2(n116), .ZN(n114) );
  NAND2_X1 U72 ( .A1(n307), .A2(n310), .ZN(n115) );
  NAND2_X1 U73 ( .A1(n308), .A2(n309), .ZN(n116) );
  NAND2_X1 U74 ( .A1(n341), .A2(n311), .ZN(n112) );
  NAND2_X1 U75 ( .A1(n92), .A2(n319), .ZN(n1) );
  OR2_X1 U76 ( .A1(n153), .A2(n152), .ZN(n130) );
  NOR2_X1 U77 ( .A1(n288), .A2(n359), .ZN(n187) );
  AND2_X1 U80 ( .A1(n2), .A2(n296), .ZN(n159) );
  AND3_X1 U81 ( .A1(n338), .A2(n295), .A3(n209), .ZN(n2) );
  INV_X1 U82 ( .A(n153), .ZN(n338) );
  NAND2_X1 U83 ( .A1(n305), .A2(n306), .ZN(n133) );
  NAND2_X1 U84 ( .A1(n352), .A2(n290), .ZN(n181) );
  NAND2_X1 U85 ( .A1(n303), .A2(n304), .ZN(n134) );
  AND2_X1 U86 ( .A1(n23), .A2(n299), .ZN(n26) );
  AND2_X1 U87 ( .A1(n144), .A2(n303), .ZN(n141) );
  NAND4_X1 U88 ( .A1(n315), .A2(n318), .A3(n317), .A4(n316), .ZN(n88) );
  NAND4_X1 U89 ( .A1(n311), .A2(n314), .A3(n313), .A4(n312), .ZN(n87) );
  NOR2_X1 U90 ( .A1(n81), .A2(n82), .ZN(n80) );
  NAND2_X1 U92 ( .A1(n319), .A2(n321), .ZN(n82) );
  NAND2_X1 U93 ( .A1(n322), .A2(n323), .ZN(n81) );
  INV_X1 U95 ( .A(n34), .ZN(n353) );
  NAND2_X1 U96 ( .A1(n182), .A2(n183), .ZN(n152) );
  NOR2_X1 U100 ( .A1(n178), .A2(n179), .ZN(n182) );
  NOR2_X1 U101 ( .A1(B[15]), .A2(n177), .ZN(n183) );
  AND2_X1 U102 ( .A1(n203), .A2(n204), .ZN(n209) );
  NOR2_X1 U103 ( .A1(n178), .A2(n179), .ZN(n203) );
  NOR2_X1 U104 ( .A1(B[15]), .A2(n177), .ZN(n204) );
  NAND2_X1 U105 ( .A1(n31), .A2(n289), .ZN(n177) );
  NOR2_X1 U106 ( .A1(n353), .A2(n359), .ZN(n10) );
  NOR2_X1 U107 ( .A1(n179), .A2(n356), .ZN(n34) );
  INV_X1 U108 ( .A(n179), .ZN(n352) );
  INV_X1 U109 ( .A(n31), .ZN(n356) );
  AND2_X1 U110 ( .A1(n29), .A2(n357), .ZN(n38) );
  INV_X1 U111 ( .A(n30), .ZN(n359) );
  AND2_X1 U112 ( .A1(n352), .A2(n355), .ZN(n29) );
  NAND2_X1 U113 ( .A1(n362), .A2(n361), .ZN(n189) );
  NOR2_X1 U114 ( .A1(n192), .A2(n193), .ZN(n9) );
  NAND2_X1 U115 ( .A1(n352), .A2(n30), .ZN(n193) );
  NOR2_X1 U116 ( .A1(n356), .A2(n189), .ZN(n188) );
  XNOR2_X1 U117 ( .A(n152), .B(n290), .ZN(DIFF[16]) );
  XNOR2_X1 U119 ( .A(n27), .B(n291), .ZN(DIFF[17]) );
  AND2_X1 U120 ( .A1(n7), .A2(n8), .ZN(n27) );
  NOR2_X1 U121 ( .A1(n178), .A2(n181), .ZN(n7) );
  XNOR2_X1 U122 ( .A(n295), .B(n130), .ZN(DIFF[20]) );
  XNOR2_X1 U123 ( .A(n302), .B(n150), .ZN(DIFF[27]) );
  NAND2_X1 U124 ( .A1(n301), .A2(n151), .ZN(n150) );
  XNOR2_X1 U125 ( .A(n298), .B(n158), .ZN(DIFF[23]) );
  NAND2_X1 U126 ( .A1(n297), .A2(n159), .ZN(n158) );
  XNOR2_X1 U127 ( .A(n139), .B(n306), .ZN(DIFF[31]) );
  NAND2_X1 U128 ( .A1(n140), .A2(n305), .ZN(n139) );
  XNOR2_X1 U129 ( .A(n310), .B(n121), .ZN(DIFF[35]) );
  NAND2_X1 U130 ( .A1(n309), .A2(n122), .ZN(n121) );
  XNOR2_X1 U131 ( .A(n110), .B(B[38]), .ZN(DIFF[38]) );
  XNOR2_X1 U132 ( .A(n318), .B(n97), .ZN(DIFF[43]) );
  NAND2_X1 U136 ( .A1(n317), .A2(n98), .ZN(n97) );
  XNOR2_X1 U137 ( .A(n323), .B(n89), .ZN(DIFF[47]) );
  NAND2_X1 U138 ( .A1(n322), .A2(n90), .ZN(n89) );
  XNOR2_X1 U148 ( .A(n208), .B(n314), .ZN(DIFF[39]) );
  NAND2_X1 U149 ( .A1(n313), .A2(n110), .ZN(n208) );
  XNOR2_X1 U150 ( .A(n327), .B(n72), .ZN(DIFF[51]) );
  NAND2_X1 U151 ( .A1(n326), .A2(n17), .ZN(n72) );
  XNOR2_X1 U152 ( .A(n331), .B(n63), .ZN(DIFF[55]) );
  NAND2_X1 U153 ( .A1(n330), .A2(n18), .ZN(n63) );
  XNOR2_X1 U154 ( .A(n335), .B(n54), .ZN(DIFF[59]) );
  NAND2_X1 U155 ( .A1(n334), .A2(n19), .ZN(n54) );
  NAND2_X1 U156 ( .A1(n41), .A2(n337), .ZN(n207) );
  NAND2_X1 U157 ( .A1(n360), .A2(n199), .ZN(n16) );
  NAND2_X1 U158 ( .A1(n358), .A2(n38), .ZN(n205) );
  NOR2_X1 U159 ( .A1(n28), .A2(B[9]), .ZN(n199) );
  NAND2_X1 U160 ( .A1(n200), .A2(n201), .ZN(n179) );
  NOR2_X1 U161 ( .A1(B[1]), .A2(\B[0] ), .ZN(n200) );
  NOR2_X1 U162 ( .A1(B[3]), .A2(B[2]), .ZN(n201) );
  AND2_X1 U163 ( .A1(n12), .A2(n13), .ZN(n30) );
  NOR2_X1 U164 ( .A1(B[11]), .A2(B[10]), .ZN(n12) );
  NOR2_X1 U165 ( .A1(B[9]), .A2(B[8]), .ZN(n13) );
  AND2_X1 U166 ( .A1(n14), .A2(n15), .ZN(n31) );
  NOR2_X1 U167 ( .A1(B[5]), .A2(B[4]), .ZN(n14) );
  NOR2_X1 U168 ( .A1(B[7]), .A2(B[6]), .ZN(n15) );
  XNOR2_X1 U169 ( .A(B[8]), .B(n34), .ZN(DIFF[8]) );
  XNOR2_X1 U170 ( .A(B[2]), .B(n32), .ZN(DIFF[2]) );
  XNOR2_X1 U171 ( .A(B[3]), .B(n206), .ZN(DIFF[3]) );
  NOR2_X1 U172 ( .A1(n350), .A2(B[2]), .ZN(n206) );
  INV_X1 U173 ( .A(n32), .ZN(n350) );
  NAND2_X1 U174 ( .A1(n184), .A2(n30), .ZN(n178) );
  NOR2_X1 U175 ( .A1(B[13]), .A2(B[12]), .ZN(n184) );
  XNOR2_X1 U176 ( .A(n362), .B(n195), .ZN(DIFF[13]) );
  NAND4_X1 U177 ( .A1(n352), .A2(n30), .A3(n196), .A4(n31), .ZN(n195) );
  NOR2_X1 U178 ( .A1(B[1]), .A2(B[12]), .ZN(n196) );
  OR2_X1 U179 ( .A1(B[8]), .A2(n353), .ZN(n28) );
  INV_X1 U180 ( .A(B[13]), .ZN(n362) );
  AND2_X1 U181 ( .A1(n354), .A2(n351), .ZN(n32) );
  INV_X1 U182 ( .A(\B[0] ), .ZN(n351) );
  INV_X1 U183 ( .A(B[12]), .ZN(n361) );
  INV_X1 U184 ( .A(B[1]), .ZN(n354) );
  INV_X1 U185 ( .A(B[6]), .ZN(n358) );
  INV_X1 U186 ( .A(B[10]), .ZN(n360) );
  INV_X1 U187 ( .A(B[4]), .ZN(n355) );
  INV_X1 U188 ( .A(B[5]), .ZN(n357) );
  XNOR2_X1 U189 ( .A(n354), .B(\B[0] ), .ZN(DIFF[1]) );
  INV_X1 U190 ( .A(n289), .ZN(n288) );
  INV_X1 U191 ( .A(B[16]), .ZN(n290) );
  INV_X1 U192 ( .A(n292), .ZN(n291) );
  INV_X1 U193 ( .A(B[17]), .ZN(n292) );
  INV_X1 U194 ( .A(B[18]), .ZN(n293) );
  INV_X1 U195 ( .A(B[19]), .ZN(n294) );
  INV_X1 U196 ( .A(B[20]), .ZN(n295) );
  INV_X1 U197 ( .A(B[21]), .ZN(n296) );
  INV_X1 U198 ( .A(B[22]), .ZN(n297) );
  INV_X1 U199 ( .A(B[23]), .ZN(n298) );
  INV_X1 U200 ( .A(B[24]), .ZN(n299) );
  INV_X1 U201 ( .A(B[25]), .ZN(n300) );
  INV_X1 U202 ( .A(B[26]), .ZN(n301) );
  INV_X1 U203 ( .A(B[27]), .ZN(n302) );
  INV_X1 U204 ( .A(B[28]), .ZN(n303) );
  INV_X1 U205 ( .A(B[29]), .ZN(n304) );
  INV_X1 U209 ( .A(B[30]), .ZN(n305) );
  INV_X1 U210 ( .A(B[31]), .ZN(n306) );
  INV_X1 U212 ( .A(B[32]), .ZN(n307) );
  INV_X1 U214 ( .A(B[33]), .ZN(n308) );
  INV_X1 U215 ( .A(B[34]), .ZN(n309) );
  INV_X1 U216 ( .A(B[35]), .ZN(n310) );
  INV_X1 U217 ( .A(B[36]), .ZN(n311) );
  INV_X1 U218 ( .A(B[37]), .ZN(n312) );
  INV_X1 U219 ( .A(B[38]), .ZN(n313) );
  INV_X1 U220 ( .A(B[39]), .ZN(n314) );
  INV_X1 U221 ( .A(B[40]), .ZN(n315) );
  INV_X1 U222 ( .A(B[41]), .ZN(n316) );
  INV_X1 U223 ( .A(B[42]), .ZN(n317) );
  INV_X1 U224 ( .A(B[43]), .ZN(n318) );
  INV_X1 U225 ( .A(B[44]), .ZN(n319) );
  INV_X1 U226 ( .A(n321), .ZN(n320) );
  INV_X1 U227 ( .A(B[45]), .ZN(n321) );
  INV_X1 U228 ( .A(B[46]), .ZN(n322) );
  INV_X1 U229 ( .A(B[47]), .ZN(n323) );
  INV_X1 U230 ( .A(B[48]), .ZN(n324) );
  INV_X1 U231 ( .A(B[49]), .ZN(n325) );
  INV_X1 U232 ( .A(B[50]), .ZN(n326) );
  INV_X1 U233 ( .A(B[51]), .ZN(n327) );
  INV_X1 U234 ( .A(B[52]), .ZN(n328) );
  INV_X1 U235 ( .A(B[53]), .ZN(n329) );
  INV_X1 U236 ( .A(B[54]), .ZN(n330) );
  INV_X1 U237 ( .A(B[55]), .ZN(n331) );
  INV_X1 U242 ( .A(B[56]), .ZN(n332) );
  INV_X1 U243 ( .A(B[57]), .ZN(n333) );
  INV_X1 U244 ( .A(B[58]), .ZN(n334) );
  INV_X1 U245 ( .A(B[59]), .ZN(n335) );
  INV_X1 U246 ( .A(B[60]), .ZN(n336) );
  INV_X1 U247 ( .A(B[62]), .ZN(n337) );
endmodule


module complement_NBIT64_18 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_18_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_17_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n5, n6, n7, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n41, n43, n44, n45, n47, n49, n51,
         n52, n58, n61, n64, n65, n70, n73, n76, n77, n82, n85, n88, n89, n91,
         n92, n93, n96, n98, n99, n101, n102, n105, n106, n114, n116, n117,
         n119, n120, n121, n122, n125, n126, n127, n131, n132, n135, n136,
         n137, n142, n143, n144, n147, n152, n153, n155, n156, n160, n166,
         n170, n171, n172, n173, n174, n178, n180, n181, n182, n183, n184,
         n186, n187, n188, n190, n191, n192, n194, n195, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U10 ( .A(n6), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U12 ( .A(n7), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U16 ( .A(n9), .B(B[12]), .Z(DIFF[12]) );
  XOR2_X1 U22 ( .A(n12), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U42 ( .A(n311), .B(n327), .Z(DIFF[49]) );
  XOR2_X1 U43 ( .A(n315), .B(n328), .Z(DIFF[53]) );
  XOR2_X1 U47 ( .A(n82), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U50 ( .A(B[47]), .B(n98), .Z(DIFF[47]) );
  XOR2_X1 U52 ( .A(n70), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U54 ( .A(n319), .B(n329), .Z(DIFF[57]) );
  XOR2_X1 U55 ( .A(n58), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U75 ( .A(n117), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U76 ( .A(n14), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U81 ( .A(n102), .B(B[40]), .Z(DIFF[40]) );
  XOR2_X1 U86 ( .A(n2), .B(n306), .Z(DIFF[45]) );
  XOR2_X1 U88 ( .A(n325), .B(B[32]), .Z(DIFF[32]) );
  XOR2_X1 U96 ( .A(n290), .B(n19), .Z(DIFF[29]) );
  XOR2_X1 U97 ( .A(n287), .B(n17), .Z(DIFF[26]) );
  XOR2_X1 U103 ( .A(n286), .B(n153), .Z(DIFF[25]) );
  XOR2_X1 U112 ( .A(n291), .B(n16), .Z(DIFF[30]) );
  XOR2_X1 U113 ( .A(n289), .B(n147), .Z(DIFF[28]) );
  XOR2_X1 U114 ( .A(n282), .B(n3), .Z(DIFF[21]) );
  XOR2_X1 U115 ( .A(n283), .B(n18), .Z(DIFF[22]) );
  XOR2_X1 U116 ( .A(n285), .B(n5), .Z(DIFF[24]) );
  XOR2_X1 U117 ( .A(n277), .B(n1), .Z(DIFF[16]) );
  XOR2_X1 U129 ( .A(n297), .B(n326), .Z(DIFF[36]) );
  XOR2_X1 U151 ( .A(B[27]), .B(n152), .Z(DIFF[27]) );
  XOR2_X1 U154 ( .A(B[23]), .B(n160), .Z(DIFF[23]) );
  XOR2_X1 U156 ( .A(B[35]), .B(n125), .Z(DIFF[35]) );
  XOR2_X1 U159 ( .A(B[43]), .B(n105), .Z(DIFF[43]) );
  XOR2_X1 U179 ( .A(n339), .B(n22), .Z(DIFF[2]) );
  XOR2_X1 U180 ( .A(n44), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U181 ( .A(n21), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U182 ( .A(n336), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U190 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U193 ( .A(B[7]), .B(n41), .Z(DIFF[7]) );
  XOR2_X1 U196 ( .A(B[14]), .B(n182), .Z(DIFF[14]) );
  NAND3_X1 U229 ( .A1(n320), .A2(n321), .A3(n319), .ZN(n52) );
  NAND3_X1 U231 ( .A1(n316), .A2(n317), .A3(n315), .ZN(n65) );
  NAND3_X1 U233 ( .A1(n312), .A2(n313), .A3(n311), .ZN(n77) );
  NAND3_X1 U235 ( .A1(n334), .A2(n20), .A3(n91), .ZN(n89) );
  NAND3_X1 U243 ( .A1(n333), .A2(n332), .A3(n135), .ZN(n132) );
  XOR2_X1 U3 ( .A(n190), .B(n313), .Z(DIFF[51]) );
  XOR2_X1 U6 ( .A(n191), .B(n317), .Z(DIFF[55]) );
  XOR2_X1 U8 ( .A(n192), .B(n321), .Z(DIFF[59]) );
  XOR2_X1 U36 ( .A(n61), .B(n318), .Z(DIFF[56]) );
  XOR2_X1 U38 ( .A(n85), .B(n310), .Z(DIFF[48]) );
  XOR2_X1 U39 ( .A(n73), .B(n314), .Z(DIFF[52]) );
  XOR2_X1 U40 ( .A(n323), .B(n47), .Z(DIFF[61]) );
  XOR2_X1 U41 ( .A(n45), .B(n324), .Z(DIFF[62]) );
  XOR2_X1 U44 ( .A(n322), .B(n49), .Z(DIFF[60]) );
  XOR2_X1 U45 ( .A(n194), .B(B[63]), .Z(DIFF[63]) );
  INV_X1 U4 ( .A(n64), .ZN(n328) );
  INV_X1 U5 ( .A(n51), .ZN(n329) );
  NOR2_X1 U7 ( .A1(n82), .A2(B[50]), .ZN(n190) );
  NOR2_X1 U9 ( .A1(n70), .A2(B[54]), .ZN(n191) );
  NOR2_X1 U11 ( .A1(n58), .A2(B[58]), .ZN(n192) );
  NOR2_X1 U13 ( .A1(n64), .A2(n65), .ZN(n61) );
  NOR2_X1 U14 ( .A1(n51), .A2(n52), .ZN(n49) );
  NAND2_X1 U15 ( .A1(n73), .A2(n314), .ZN(n64) );
  NAND2_X1 U17 ( .A1(n61), .A2(n318), .ZN(n51) );
  NAND2_X1 U18 ( .A1(n311), .A2(n327), .ZN(n82) );
  NAND2_X1 U19 ( .A1(n315), .A2(n328), .ZN(n70) );
  NAND2_X1 U20 ( .A1(n319), .A2(n329), .ZN(n58) );
  AND2_X1 U21 ( .A1(n323), .A2(n47), .ZN(n45) );
  AND2_X1 U23 ( .A1(n322), .A2(n49), .ZN(n47) );
  NOR2_X1 U24 ( .A1(B[32]), .A2(n325), .ZN(n127) );
  NAND2_X1 U25 ( .A1(n308), .A2(n99), .ZN(n98) );
  NOR2_X1 U26 ( .A1(n76), .A2(n77), .ZN(n73) );
  XNOR2_X1 U27 ( .A(n99), .B(B[46]), .ZN(DIFF[46]) );
  INV_X1 U28 ( .A(n76), .ZN(n327) );
  NAND2_X1 U29 ( .A1(n308), .A2(n309), .ZN(n92) );
  NAND2_X1 U30 ( .A1(n45), .A2(n324), .ZN(n194) );
  NOR2_X1 U31 ( .A1(n117), .A2(B[37]), .ZN(n116) );
  NOR2_X1 U32 ( .A1(n2), .A2(n306), .ZN(n99) );
  NOR2_X1 U33 ( .A1(n14), .A2(B[41]), .ZN(n106) );
  NAND2_X1 U34 ( .A1(n20), .A2(n326), .ZN(n102) );
  INV_X1 U35 ( .A(n88), .ZN(n326) );
  NAND2_X1 U37 ( .A1(n101), .A2(n305), .ZN(n2) );
  NAND2_X1 U46 ( .A1(n326), .A2(n297), .ZN(n117) );
  OR2_X1 U48 ( .A1(B[40]), .A2(n102), .ZN(n14) );
  INV_X1 U49 ( .A(n119), .ZN(n325) );
  NAND2_X1 U51 ( .A1(n85), .A2(n310), .ZN(n76) );
  NOR2_X1 U53 ( .A1(n102), .A2(n96), .ZN(n101) );
  NOR2_X1 U56 ( .A1(n131), .A2(n132), .ZN(n119) );
  NOR2_X1 U57 ( .A1(n136), .A2(n137), .ZN(n135) );
  INV_X1 U58 ( .A(n143), .ZN(n333) );
  NOR2_X1 U59 ( .A1(n331), .A2(n143), .ZN(n147) );
  XNOR2_X1 U60 ( .A(n126), .B(B[34]), .ZN(DIFF[34]) );
  XNOR2_X1 U61 ( .A(n281), .B(n131), .ZN(DIFF[20]) );
  XOR2_X1 U62 ( .A(n276), .B(B[18]), .Z(DIFF[18]) );
  NAND2_X1 U63 ( .A1(n15), .A2(n278), .ZN(n276) );
  XNOR2_X1 U64 ( .A(n15), .B(B[17]), .ZN(DIFF[17]) );
  NAND2_X1 U65 ( .A1(n119), .A2(n120), .ZN(n88) );
  NOR2_X1 U66 ( .A1(n121), .A2(n122), .ZN(n120) );
  NAND2_X1 U67 ( .A1(n294), .A2(n295), .ZN(n122) );
  NAND2_X1 U68 ( .A1(n293), .A2(n296), .ZN(n121) );
  AND2_X1 U69 ( .A1(n127), .A2(n294), .ZN(n126) );
  INV_X1 U70 ( .A(B[17]), .ZN(n278) );
  AND2_X1 U71 ( .A1(n153), .A2(n286), .ZN(n17) );
  AND2_X1 U72 ( .A1(n3), .A2(n282), .ZN(n18) );
  INV_X1 U73 ( .A(n156), .ZN(n330) );
  NAND2_X1 U74 ( .A1(n291), .A2(n292), .ZN(n136) );
  XNOR2_X1 U77 ( .A(n144), .B(n292), .ZN(DIFF[31]) );
  NAND2_X1 U78 ( .A1(n16), .A2(n291), .ZN(n144) );
  AND2_X1 U79 ( .A1(n19), .A2(n290), .ZN(n16) );
  XNOR2_X1 U80 ( .A(n300), .B(n195), .ZN(DIFF[39]) );
  NAND2_X1 U82 ( .A1(n299), .A2(n116), .ZN(n195) );
  NAND2_X1 U83 ( .A1(n289), .A2(n290), .ZN(n137) );
  INV_X1 U84 ( .A(n5), .ZN(n331) );
  AND2_X1 U85 ( .A1(n147), .A2(n289), .ZN(n19) );
  NAND2_X1 U87 ( .A1(n295), .A2(n126), .ZN(n125) );
  INV_X1 U89 ( .A(n142), .ZN(n332) );
  NOR2_X1 U90 ( .A1(n88), .A2(n89), .ZN(n85) );
  INV_X1 U91 ( .A(n96), .ZN(n334) );
  NOR2_X1 U92 ( .A1(n92), .A2(n93), .ZN(n91) );
  XNOR2_X1 U93 ( .A(B[44]), .B(n101), .ZN(DIFF[44]) );
  AND4_X1 U94 ( .A1(n297), .A2(n300), .A3(n299), .A4(n298), .ZN(n20) );
  NAND2_X1 U95 ( .A1(n305), .A2(n307), .ZN(n93) );
  INV_X1 U98 ( .A(n173), .ZN(n335) );
  INV_X1 U99 ( .A(n184), .ZN(n336) );
  NAND2_X1 U100 ( .A1(n166), .A2(n1), .ZN(n6) );
  NAND2_X1 U101 ( .A1(n303), .A2(n106), .ZN(n105) );
  NAND2_X1 U102 ( .A1(n287), .A2(n17), .ZN(n152) );
  NAND2_X1 U104 ( .A1(n178), .A2(n342), .ZN(n7) );
  INV_X1 U105 ( .A(n180), .ZN(n342) );
  NOR2_X1 U106 ( .A1(n173), .A2(n181), .ZN(n178) );
  NAND4_X1 U107 ( .A1(n281), .A2(n284), .A3(n283), .A4(n282), .ZN(n142) );
  NAND4_X1 U108 ( .A1(n277), .A2(n280), .A3(n279), .A4(n278), .ZN(n156) );
  NAND4_X1 U109 ( .A1(n285), .A2(n288), .A3(n287), .A4(n286), .ZN(n143) );
  XNOR2_X1 U110 ( .A(B[33]), .B(n127), .ZN(DIFF[33]) );
  NOR2_X1 U111 ( .A1(B[24]), .A2(n331), .ZN(n153) );
  XNOR2_X1 U118 ( .A(n116), .B(B[38]), .ZN(DIFF[38]) );
  XNOR2_X1 U119 ( .A(n106), .B(B[42]), .ZN(DIFF[42]) );
  NAND2_X1 U120 ( .A1(n330), .A2(n1), .ZN(n131) );
  AND3_X1 U121 ( .A1(n281), .A2(n330), .A3(n1), .ZN(n3) );
  AND2_X1 U122 ( .A1(n1), .A2(n277), .ZN(n15) );
  AND2_X1 U123 ( .A1(n155), .A2(n1), .ZN(n5) );
  NOR2_X1 U124 ( .A1(n142), .A2(n156), .ZN(n155) );
  NAND2_X1 U125 ( .A1(n283), .A2(n18), .ZN(n160) );
  NAND4_X1 U126 ( .A1(n301), .A2(n304), .A3(n303), .A4(n302), .ZN(n96) );
  NOR2_X1 U127 ( .A1(n173), .A2(n180), .ZN(n183) );
  NOR2_X1 U128 ( .A1(n173), .A2(n172), .ZN(n184) );
  NAND2_X1 U130 ( .A1(n335), .A2(n341), .ZN(n44) );
  INV_X1 U131 ( .A(n24), .ZN(n344) );
  NAND4_X1 U132 ( .A1(n338), .A2(n337), .A3(n339), .A4(n340), .ZN(n173) );
  AND2_X1 U133 ( .A1(n338), .A2(n337), .ZN(n22) );
  NAND2_X1 U134 ( .A1(n346), .A2(n347), .ZN(n181) );
  AND3_X1 U135 ( .A1(n170), .A2(n335), .A3(n171), .ZN(n1) );
  NOR3_X1 U136 ( .A1(n174), .A2(B[12]), .A3(n344), .ZN(n170) );
  NOR2_X1 U137 ( .A1(B[15]), .A2(n172), .ZN(n171) );
  NAND2_X1 U138 ( .A1(n346), .A2(n347), .ZN(n174) );
  NOR2_X1 U139 ( .A1(n44), .A2(B[5]), .ZN(n43) );
  NOR2_X1 U140 ( .A1(n21), .A2(B[9]), .ZN(n186) );
  NAND2_X1 U141 ( .A1(n346), .A2(n183), .ZN(n182) );
  NAND2_X1 U142 ( .A1(n24), .A2(n184), .ZN(n9) );
  NAND2_X1 U143 ( .A1(n343), .A2(n43), .ZN(n41) );
  INV_X1 U144 ( .A(B[6]), .ZN(n343) );
  NAND2_X1 U145 ( .A1(n345), .A2(n186), .ZN(n12) );
  INV_X1 U146 ( .A(B[10]), .ZN(n345) );
  XNOR2_X1 U147 ( .A(n183), .B(B[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U148 ( .A(n43), .B(B[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U149 ( .A(n186), .B(B[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U150 ( .A(n173), .B(n341), .ZN(DIFF[4]) );
  XNOR2_X1 U152 ( .A(n114), .B(n340), .ZN(DIFF[3]) );
  NAND2_X1 U153 ( .A1(n22), .A2(n339), .ZN(n114) );
  NAND2_X1 U155 ( .A1(n187), .A2(n188), .ZN(n172) );
  NOR2_X1 U157 ( .A1(B[5]), .A2(B[4]), .ZN(n187) );
  NOR2_X1 U158 ( .A1(B[6]), .A2(B[7]), .ZN(n188) );
  AND2_X1 U160 ( .A1(n10), .A2(n11), .ZN(n24) );
  NOR2_X1 U161 ( .A1(B[11]), .A2(B[10]), .ZN(n10) );
  NOR2_X1 U162 ( .A1(B[9]), .A2(B[8]), .ZN(n11) );
  OR2_X1 U163 ( .A1(n23), .A2(n172), .ZN(n180) );
  OR2_X1 U164 ( .A1(B[12]), .A2(n344), .ZN(n23) );
  OR2_X1 U165 ( .A1(B[8]), .A2(n336), .ZN(n21) );
  INV_X1 U166 ( .A(B[13]), .ZN(n346) );
  INV_X1 U167 ( .A(B[2]), .ZN(n339) );
  INV_X1 U168 ( .A(B[3]), .ZN(n340) );
  INV_X1 U169 ( .A(B[4]), .ZN(n341) );
  INV_X1 U170 ( .A(B[14]), .ZN(n347) );
  INV_X1 U171 ( .A(\B[0] ), .ZN(n337) );
  INV_X1 U172 ( .A(B[1]), .ZN(n338) );
  NOR3_X1 U173 ( .A1(B[16]), .A2(B[17]), .A3(B[18]), .ZN(n166) );
  INV_X1 U174 ( .A(B[16]), .ZN(n277) );
  INV_X1 U175 ( .A(B[18]), .ZN(n279) );
  INV_X1 U176 ( .A(B[19]), .ZN(n280) );
  INV_X1 U177 ( .A(B[20]), .ZN(n281) );
  INV_X1 U178 ( .A(B[21]), .ZN(n282) );
  INV_X1 U183 ( .A(B[22]), .ZN(n283) );
  INV_X1 U184 ( .A(B[23]), .ZN(n284) );
  INV_X1 U185 ( .A(B[24]), .ZN(n285) );
  INV_X1 U186 ( .A(B[25]), .ZN(n286) );
  INV_X1 U187 ( .A(B[26]), .ZN(n287) );
  INV_X1 U188 ( .A(B[27]), .ZN(n288) );
  INV_X1 U189 ( .A(B[28]), .ZN(n289) );
  INV_X1 U191 ( .A(B[29]), .ZN(n290) );
  INV_X1 U192 ( .A(B[30]), .ZN(n291) );
  INV_X1 U194 ( .A(B[31]), .ZN(n292) );
  INV_X1 U195 ( .A(B[32]), .ZN(n293) );
  INV_X1 U197 ( .A(B[33]), .ZN(n294) );
  INV_X1 U198 ( .A(B[34]), .ZN(n295) );
  INV_X1 U199 ( .A(B[35]), .ZN(n296) );
  INV_X1 U200 ( .A(B[36]), .ZN(n297) );
  INV_X1 U201 ( .A(B[37]), .ZN(n298) );
  INV_X1 U202 ( .A(B[38]), .ZN(n299) );
  INV_X1 U203 ( .A(B[39]), .ZN(n300) );
  INV_X1 U204 ( .A(B[40]), .ZN(n301) );
  INV_X1 U205 ( .A(B[41]), .ZN(n302) );
  INV_X1 U206 ( .A(B[42]), .ZN(n303) );
  INV_X1 U207 ( .A(B[43]), .ZN(n304) );
  INV_X1 U208 ( .A(B[44]), .ZN(n305) );
  INV_X1 U209 ( .A(n307), .ZN(n306) );
  INV_X1 U210 ( .A(B[45]), .ZN(n307) );
  INV_X1 U211 ( .A(B[46]), .ZN(n308) );
  INV_X1 U212 ( .A(B[47]), .ZN(n309) );
  INV_X1 U213 ( .A(B[48]), .ZN(n310) );
  INV_X1 U214 ( .A(B[49]), .ZN(n311) );
  INV_X1 U215 ( .A(B[50]), .ZN(n312) );
  INV_X1 U216 ( .A(B[51]), .ZN(n313) );
  INV_X1 U217 ( .A(B[52]), .ZN(n314) );
  INV_X1 U218 ( .A(B[53]), .ZN(n315) );
  INV_X1 U219 ( .A(B[54]), .ZN(n316) );
  INV_X1 U220 ( .A(B[55]), .ZN(n317) );
  INV_X1 U221 ( .A(B[56]), .ZN(n318) );
  INV_X1 U222 ( .A(B[57]), .ZN(n319) );
  INV_X1 U223 ( .A(B[58]), .ZN(n320) );
  INV_X1 U224 ( .A(B[59]), .ZN(n321) );
  INV_X1 U225 ( .A(B[60]), .ZN(n322) );
  INV_X1 U226 ( .A(B[61]), .ZN(n323) );
  INV_X1 U227 ( .A(B[62]), .ZN(n324) );
endmodule


module complement_NBIT64_17 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_17_DW01_sub_2 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_16_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U2 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U4 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U5 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U6 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U7 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U8 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U9 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U10 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U11 ( .A(n205), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U12 ( .A1(n243), .A2(B[17]), .ZN(n205) );
  OR3_X1 U13 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U14 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U15 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U16 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U17 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U18 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U19 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U20 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U21 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U22 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U23 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U24 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U25 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U26 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U27 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U28 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U29 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U30 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U31 ( .A(n231), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U32 ( .A1(n239), .A2(B[21]), .ZN(n231) );
  XNOR2_X1 U33 ( .A(n227), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U34 ( .A1(n235), .A2(B[25]), .ZN(n227) );
  XNOR2_X1 U35 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U36 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U37 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U38 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U39 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U40 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  XNOR2_X1 U41 ( .A(n209), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U42 ( .A1(n226), .A2(B[33]), .ZN(n209) );
  XNOR2_X1 U43 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U44 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U45 ( .A(n236), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U46 ( .A1(n222), .A2(B[37]), .ZN(n236) );
  XNOR2_X1 U47 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U48 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U49 ( .A(n215), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U50 ( .A1(n218), .A2(B[41]), .ZN(n215) );
  XNOR2_X1 U51 ( .A(n219), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U52 ( .A1(n214), .A2(B[45]), .ZN(n219) );
  XNOR2_X1 U53 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U54 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U55 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U56 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U57 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U58 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U59 ( .A(n193), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U60 ( .A1(n204), .A2(B[53]), .ZN(n193) );
  XNOR2_X1 U61 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U62 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U63 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U64 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U65 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U66 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U67 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U68 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U69 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U70 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U71 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U72 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  OR3_X1 U73 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U74 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U75 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U76 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U77 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U78 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U79 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U80 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U83 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U84 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U88 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U91 ( .A(n240), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U94 ( .A1(n190), .A2(B[9]), .ZN(n240) );
  XNOR2_X1 U97 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U100 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  OR3_X1 U104 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U107 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U110 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U113 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U116 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_16 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_16_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_15_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U3 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U5 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U6 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U7 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U8 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U9 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U10 ( .A(n193), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U11 ( .A1(n204), .A2(B[53]), .ZN(n193) );
  XNOR2_X1 U12 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U13 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  OR3_X1 U14 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U15 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U16 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U17 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U18 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U20 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U21 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U22 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U23 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U24 ( .A(n205), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U25 ( .A1(n222), .A2(B[37]), .ZN(n205) );
  OR3_X1 U26 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U27 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U28 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  XNOR2_X1 U29 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U30 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U31 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U32 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U33 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U34 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U35 ( .A(n236), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U36 ( .A1(n230), .A2(B[29]), .ZN(n236) );
  XNOR2_X1 U37 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U38 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U39 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U40 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U41 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U42 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U43 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U44 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  XNOR2_X1 U45 ( .A(n209), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U46 ( .A1(n239), .A2(B[21]), .ZN(n209) );
  XNOR2_X1 U47 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U48 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U49 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U50 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U51 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U52 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U53 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U54 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  NOR2_X1 U55 ( .A1(n243), .A2(B[17]), .ZN(n223) );
  OR3_X1 U56 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U57 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U58 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U59 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U60 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U61 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U62 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U63 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U64 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U65 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U66 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U67 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U68 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U69 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U70 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U71 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U72 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U73 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U74 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U75 ( .A(n240), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U76 ( .A1(n194), .A2(B[5]), .ZN(n240) );
  XNOR2_X1 U77 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U78 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U79 ( .A(n248), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U80 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  XNOR2_X1 U83 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U84 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U88 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U91 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U94 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U97 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U100 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U104 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U107 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(n223), .B(B[18]), .ZN(DIFF[18]) );
  OR3_X1 U123 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_15 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_15_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_14_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U6 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U3 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U4 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U5 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U7 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U8 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U9 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U10 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U11 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U12 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U13 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U14 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U15 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U16 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U17 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U18 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U19 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U20 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U21 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U22 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U23 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U24 ( .A(n205), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U25 ( .A1(n239), .A2(B[21]), .ZN(n205) );
  XNOR2_X1 U26 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U27 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U28 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U29 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U30 ( .A(n236), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U31 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  XNOR2_X1 U32 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U33 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  XNOR2_X1 U34 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U35 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U36 ( .A(n215), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U37 ( .A1(n222), .A2(B[37]), .ZN(n215) );
  XNOR2_X1 U38 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U39 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U40 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U41 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U42 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U43 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U44 ( .A(n223), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U45 ( .A1(n214), .A2(B[45]), .ZN(n223) );
  XNOR2_X1 U46 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U47 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR2_X1 U48 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  XNOR2_X1 U49 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U50 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U51 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U52 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U53 ( .A(n189), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U54 ( .A1(n243), .A2(B[17]), .ZN(n189) );
  XNOR2_X1 U55 ( .A(n193), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U56 ( .A1(n196), .A2(B[62]), .ZN(n193) );
  XNOR2_X1 U57 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U58 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U59 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U60 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U61 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U62 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U63 ( .A(n201), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U64 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  XNOR2_X1 U65 ( .A(n227), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U66 ( .A1(n218), .A2(B[41]), .ZN(n227) );
  XNOR2_X1 U67 ( .A(n231), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U68 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR3_X1 U69 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  XNOR2_X1 U70 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U71 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U72 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U73 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U74 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U75 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U76 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U77 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U78 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U79 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U80 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U83 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U84 ( .A(n240), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U88 ( .A1(n190), .A2(B[9]), .ZN(n240) );
  XNOR2_X1 U91 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U97 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  OR3_X1 U100 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U104 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U107 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U110 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U113 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U116 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_14 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_14_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_13_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n215, n219,
         n223, n227, n231, n236, n240, n244, n248, n252, n253;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U5 ( .A(n197), .B(n253), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n253), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U3 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U4 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U8 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U9 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U10 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U11 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  OR3_X1 U12 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U13 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U14 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U15 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  OR3_X1 U16 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  XNOR2_X1 U17 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U18 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U19 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U20 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U21 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U22 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U23 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U24 ( .A(n201), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U25 ( .A1(n239), .A2(B[21]), .ZN(n201) );
  XNOR2_X1 U26 ( .A(n252), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U27 ( .A1(n208), .A2(B[49]), .ZN(n252) );
  XNOR2_X1 U28 ( .A(n231), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U29 ( .A1(n226), .A2(B[33]), .ZN(n231) );
  XNOR2_X1 U30 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U31 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U32 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U33 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U34 ( .A(n223), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U35 ( .A1(n214), .A2(B[45]), .ZN(n223) );
  XNOR2_X1 U36 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U37 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U38 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U39 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U40 ( .A(n215), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U41 ( .A1(n222), .A2(B[37]), .ZN(n215) );
  XNOR2_X1 U42 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U43 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR3_X1 U44 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U45 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U46 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U47 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U48 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U49 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U50 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U51 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U52 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U53 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U54 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U55 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U56 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  NOR2_X1 U57 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U58 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U59 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U60 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U61 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U62 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U63 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U64 ( .A(n205), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U65 ( .A1(n235), .A2(B[25]), .ZN(n205) );
  XNOR2_X1 U66 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U67 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U68 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U69 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U70 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U71 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U72 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U73 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U74 ( .A(n236), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U75 ( .A1(n194), .A2(B[5]), .ZN(n236) );
  XNOR2_X1 U76 ( .A(n240), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U77 ( .A1(n190), .A2(B[9]), .ZN(n240) );
  XNOR2_X1 U78 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U79 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  XNOR2_X1 U80 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U83 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U84 ( .A(n248), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U88 ( .A1(n243), .A2(B[17]), .ZN(n248) );
  OR3_X1 U91 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U94 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U97 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U100 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U104 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U107 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  OR3_X1 U123 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  INV_X1 U126 ( .A(B[61]), .ZN(n253) );
endmodule


module complement_NBIT64_13 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_13_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_12_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U3 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U5 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U8 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U9 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U10 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U11 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U12 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U13 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U14 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U15 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U16 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U17 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U18 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U19 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U20 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U21 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U22 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U23 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U24 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U25 ( .A(n205), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U26 ( .A1(n239), .A2(B[21]), .ZN(n205) );
  XNOR2_X1 U27 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U28 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U29 ( .A(n209), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U30 ( .A1(n222), .A2(B[37]), .ZN(n209) );
  XNOR2_X1 U31 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U32 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR2_X1 U33 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U34 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U35 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U36 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U37 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U38 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U39 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U40 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U41 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U42 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U43 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U44 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U45 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U46 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U47 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U48 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U49 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U50 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U51 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U52 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U53 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U54 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  XNOR2_X1 U55 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U56 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U57 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U58 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  XNOR2_X1 U59 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U60 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U61 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U62 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U63 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U64 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U65 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U66 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U67 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U68 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U69 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U70 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U71 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U72 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U73 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U74 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U75 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U76 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U77 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U78 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U79 ( .A(n236), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U80 ( .A1(n190), .A2(B[9]), .ZN(n236) );
  XNOR2_X1 U83 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U84 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U88 ( .A(n244), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U91 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR3_X1 U94 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U100 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U104 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U107 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U110 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U113 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U116 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_12 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_12_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_11_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n219,
         n223, n227, n231, n236, n240, n244, n248, n252, n253;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n253), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n253), .ZN(n196) );
  XNOR2_X1 U2 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U5 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U6 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  OR3_X1 U7 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  NOR3_X1 U8 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U9 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U10 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U11 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U12 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U13 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U14 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U15 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  OR3_X1 U16 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U17 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U18 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  XNOR2_X1 U19 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U20 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U21 ( .A(n201), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U22 ( .A1(n218), .A2(B[41]), .ZN(n201) );
  XNOR2_X1 U23 ( .A(n252), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U24 ( .A1(n214), .A2(B[45]), .ZN(n252) );
  XNOR2_X1 U25 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U26 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U27 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U28 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U29 ( .A(n219), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U30 ( .A1(n208), .A2(B[49]), .ZN(n219) );
  OR3_X1 U31 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U32 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U33 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U34 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U35 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U36 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U37 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U38 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U39 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U40 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U42 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U43 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  NOR2_X1 U44 ( .A1(n239), .A2(B[21]), .ZN(n209) );
  XNOR2_X1 U45 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U46 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U47 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U48 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U49 ( .A(n231), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U50 ( .A1(n226), .A2(B[33]), .ZN(n231) );
  XNOR2_X1 U51 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U52 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U53 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U54 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U55 ( .A(n223), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U56 ( .A1(n235), .A2(B[25]), .ZN(n223) );
  XNOR2_X1 U57 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U58 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U59 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U60 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U61 ( .A(n205), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U62 ( .A1(n222), .A2(B[37]), .ZN(n205) );
  XNOR2_X1 U63 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U64 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U65 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U66 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U67 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U68 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U69 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U70 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U71 ( .A(n236), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U72 ( .A1(n194), .A2(B[5]), .ZN(n236) );
  XNOR2_X1 U73 ( .A(n240), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U74 ( .A1(n190), .A2(B[9]), .ZN(n240) );
  XNOR2_X1 U75 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U76 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  XNOR2_X1 U77 ( .A(n248), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U78 ( .A1(n243), .A2(B[17]), .ZN(n248) );
  XNOR2_X1 U79 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U80 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U83 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U84 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U88 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U91 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U94 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U97 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U100 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U104 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U107 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(n209), .B(B[22]), .ZN(DIFF[22]) );
  OR3_X1 U123 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  INV_X1 U126 ( .A(B[61]), .ZN(n253) );
endmodule


module complement_NBIT64_11 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_11_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_10_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U10 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U3 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U4 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U5 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  XNOR2_X1 U7 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U8 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  XNOR2_X1 U9 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U11 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U12 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U13 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U14 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U15 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U16 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U17 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U18 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U19 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U20 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U21 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U22 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U23 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U24 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U25 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U26 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U27 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U28 ( .A(n205), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U29 ( .A1(n230), .A2(B[29]), .ZN(n205) );
  XNOR2_X1 U30 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U31 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U32 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U33 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U34 ( .A(n223), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U35 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  XNOR2_X1 U36 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U37 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U38 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U39 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U40 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U41 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U42 ( .A(n219), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U43 ( .A1(n208), .A2(B[49]), .ZN(n219) );
  XNOR2_X1 U44 ( .A(n201), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U45 ( .A1(n204), .A2(B[53]), .ZN(n201) );
  XNOR2_X1 U46 ( .A(n189), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U47 ( .A1(n239), .A2(B[21]), .ZN(n189) );
  XNOR2_X1 U48 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U49 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U50 ( .A(n195), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U51 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  XNOR2_X1 U52 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U53 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U54 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U55 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U56 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U57 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U58 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U59 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U60 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U61 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U62 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U63 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR3_X1 U64 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  XNOR2_X1 U65 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U66 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U67 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U68 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U69 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U70 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U71 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U72 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U73 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U74 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U75 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U76 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U77 ( .A(n236), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U78 ( .A1(n194), .A2(B[5]), .ZN(n236) );
  XNOR2_X1 U79 ( .A(n240), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U80 ( .A1(n190), .A2(B[9]), .ZN(n240) );
  XNOR2_X1 U83 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U84 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  XNOR2_X1 U88 ( .A(n248), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U91 ( .A1(n243), .A2(B[17]), .ZN(n248) );
  OR3_X1 U94 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U97 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U100 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U104 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U107 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U110 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U113 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U116 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_10 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_10_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_9_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U5 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U3 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U4 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U6 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U7 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U8 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U9 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  OR3_X1 U10 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  XNOR2_X1 U11 ( .A(n223), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U12 ( .A1(n235), .A2(B[25]), .ZN(n223) );
  XNOR2_X1 U13 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U14 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U15 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U16 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U17 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U19 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U20 ( .A(n227), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U21 ( .A1(n222), .A2(B[37]), .ZN(n227) );
  NOR2_X1 U22 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U23 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U24 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U25 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U26 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U27 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U28 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U29 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U30 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U31 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U32 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U33 ( .A(n195), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U34 ( .A1(n230), .A2(B[29]), .ZN(n195) );
  XNOR2_X1 U35 ( .A(n209), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U36 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  XNOR2_X1 U37 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U38 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U39 ( .A(n219), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U40 ( .A1(n204), .A2(B[53]), .ZN(n219) );
  XNOR2_X1 U41 ( .A(n215), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U42 ( .A1(n226), .A2(B[33]), .ZN(n215) );
  XNOR2_X1 U43 ( .A(n201), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U44 ( .A1(n218), .A2(B[41]), .ZN(n201) );
  XNOR2_X1 U45 ( .A(n205), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U46 ( .A1(n214), .A2(B[45]), .ZN(n205) );
  OR3_X1 U47 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U48 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U49 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U50 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U51 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U52 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U53 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U54 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U55 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U56 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U57 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U58 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U59 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U60 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U61 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U62 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U63 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U64 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U65 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U66 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U67 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U68 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U69 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U70 ( .A(n231), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U71 ( .A1(n194), .A2(B[5]), .ZN(n231) );
  XNOR2_X1 U72 ( .A(n236), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U73 ( .A1(n190), .A2(B[9]), .ZN(n236) );
  XNOR2_X1 U74 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U75 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U76 ( .A(n244), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U77 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  XNOR2_X1 U78 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U79 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U80 ( .A(n248), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U83 ( .A1(n239), .A2(B[21]), .ZN(n248) );
  OR3_X1 U84 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U88 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U91 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U94 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U97 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U100 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U104 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U107 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR3_X1 U123 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_9 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_9_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_8_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U3 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U5 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U6 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U7 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U8 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U9 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U10 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U11 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U12 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U13 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U14 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U15 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U16 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U17 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U18 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U19 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U20 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U21 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U22 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U23 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U24 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U25 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U26 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U27 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U28 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U29 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U30 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U31 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U32 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U33 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U34 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  XNOR2_X1 U35 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U36 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U37 ( .A(n223), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U38 ( .A1(n235), .A2(B[25]), .ZN(n223) );
  XNOR2_X1 U39 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U40 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U41 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U42 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U43 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U44 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U45 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U46 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U47 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U48 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U49 ( .A(n209), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U50 ( .A1(n204), .A2(B[53]), .ZN(n209) );
  XNOR2_X1 U51 ( .A(n205), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U52 ( .A1(n208), .A2(B[49]), .ZN(n205) );
  XNOR2_X1 U53 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U54 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U55 ( .A(n215), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U56 ( .A1(n222), .A2(B[37]), .ZN(n215) );
  XNOR2_X1 U57 ( .A(n195), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U58 ( .A1(n218), .A2(B[41]), .ZN(n195) );
  XNOR2_X1 U59 ( .A(n201), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U60 ( .A1(n214), .A2(B[45]), .ZN(n201) );
  OR3_X1 U61 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U62 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U63 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U64 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U65 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U66 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U67 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U68 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U69 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U70 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U71 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U72 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U73 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U74 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U75 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U76 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U77 ( .A1(n190), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U78 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U79 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U80 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U83 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U84 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U88 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  OR3_X1 U91 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U94 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U97 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U100 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U104 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U107 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U110 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U113 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U116 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_8 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_8_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_7_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  XNOR2_X1 U1 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U2 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  NAND2_X1 U3 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U5 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U8 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U9 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U10 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U11 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR3_X1 U12 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U13 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U14 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  XNOR2_X1 U15 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U16 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U17 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U18 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U19 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U20 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U21 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U22 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U23 ( .A(n209), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U24 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  XNOR2_X1 U25 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U26 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U27 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U28 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U29 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U30 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U31 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U32 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U33 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U34 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U35 ( .A(n205), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U36 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  XNOR2_X1 U37 ( .A(n201), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U38 ( .A1(n222), .A2(B[37]), .ZN(n201) );
  OR3_X1 U39 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U40 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U41 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U42 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U43 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U44 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U45 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U46 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U47 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U48 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U49 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U50 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U51 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U52 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U53 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U54 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U55 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  NOR2_X1 U56 ( .A1(n235), .A2(B[25]), .ZN(n195) );
  XNOR2_X1 U57 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U58 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U59 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U60 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U61 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U62 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U63 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U64 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U65 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U66 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U67 ( .A(n231), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U68 ( .A1(n194), .A2(B[5]), .ZN(n231) );
  XNOR2_X1 U69 ( .A(n236), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U70 ( .A1(n190), .A2(B[9]), .ZN(n236) );
  XNOR2_X1 U71 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U72 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U73 ( .A(n248), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U74 ( .A1(n239), .A2(B[21]), .ZN(n248) );
  XNOR2_X1 U75 ( .A(n244), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U76 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  XNOR2_X1 U77 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U78 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U79 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U80 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U83 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U84 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U88 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U91 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U94 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U97 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U100 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U104 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U107 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(n195), .B(B[26]), .ZN(DIFF[26]) );
  OR3_X1 U123 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_7 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_7_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_6_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n191, n192, n193, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n190, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U82 ( .A(n192), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U83 ( .A(n194), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n191), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n196), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U5 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n191) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U3 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U4 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U7 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U8 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U9 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U10 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U11 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U12 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U13 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U14 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U15 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U16 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U17 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U18 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U19 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U20 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U21 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U22 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U23 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U24 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U25 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U26 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U27 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U28 ( .A(n190), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U29 ( .A1(n191), .A2(B[62]), .ZN(n190) );
  XNOR2_X1 U30 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U31 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U32 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U33 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U34 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U35 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U36 ( .A(n209), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U37 ( .A1(n214), .A2(B[45]), .ZN(n209) );
  XNOR2_X1 U38 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U39 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U40 ( .A(n215), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U41 ( .A1(n204), .A2(B[53]), .ZN(n215) );
  OR3_X1 U42 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U43 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U44 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  XNOR2_X1 U45 ( .A(n223), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U46 ( .A1(n226), .A2(B[33]), .ZN(n223) );
  XNOR2_X1 U47 ( .A(n189), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U48 ( .A1(n235), .A2(B[25]), .ZN(n189) );
  XNOR2_X1 U49 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U50 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U51 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U52 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U53 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U54 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U55 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U56 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U57 ( .A(n205), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U58 ( .A1(n218), .A2(B[41]), .ZN(n205) );
  XNOR2_X1 U59 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U60 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U61 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U62 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U63 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U64 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U65 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U66 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U67 ( .A(B[8]), .B(n193), .ZN(DIFF[8]) );
  NOR2_X1 U68 ( .A1(B[7]), .A2(n194), .ZN(n193) );
  XNOR2_X1 U69 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U70 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U71 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U72 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U73 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U74 ( .A1(n196), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U75 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U76 ( .A1(n192), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U77 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U78 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U79 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U80 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U81 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U84 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  OR3_X1 U88 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U91 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U94 ( .A1(B[10]), .A2(B[9]), .A3(n192), .ZN(n249) );
  OR3_X1 U97 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U100 ( .A1(B[5]), .A2(B[6]), .A3(n196), .ZN(n194) );
  OR3_X1 U104 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U107 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U110 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U113 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U116 ( .A1(B[7]), .A2(B[8]), .A3(n194), .ZN(n192) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n196) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_6 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_6_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_5_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  XNOR2_X1 U1 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U2 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  NAND2_X1 U3 ( .A1(n197), .A2(n252), .ZN(n196) );
  NOR3_X1 U5 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U8 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U9 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U10 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U11 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  XNOR2_X1 U12 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U13 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U14 ( .A(n209), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U15 ( .A1(n204), .A2(B[53]), .ZN(n209) );
  XNOR2_X1 U16 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U17 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U18 ( .A(n215), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U19 ( .A1(n200), .A2(B[57]), .ZN(n215) );
  OR3_X1 U20 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U21 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U22 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U23 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U24 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U25 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U26 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U27 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U28 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U29 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U30 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U31 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U32 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  NOR2_X1 U33 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U34 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U35 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U36 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U37 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U38 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U39 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U40 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U41 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U42 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U43 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U44 ( .A(n193), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U45 ( .A1(n226), .A2(B[33]), .ZN(n193) );
  XNOR2_X1 U46 ( .A(n201), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U47 ( .A1(n218), .A2(B[41]), .ZN(n201) );
  XNOR2_X1 U48 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U49 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  XNOR2_X1 U50 ( .A(n195), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U51 ( .A1(n214), .A2(B[45]), .ZN(n195) );
  XNOR2_X1 U52 ( .A(n205), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U53 ( .A1(n208), .A2(B[49]), .ZN(n205) );
  XNOR2_X1 U54 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U55 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U56 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U57 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U58 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U59 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U60 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U61 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U62 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U63 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U64 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U65 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U66 ( .A(n227), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U67 ( .A1(n194), .A2(B[5]), .ZN(n227) );
  XNOR2_X1 U68 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U69 ( .A1(n190), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U70 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U71 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U72 ( .A(n248), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U73 ( .A1(n239), .A2(B[21]), .ZN(n248) );
  XNOR2_X1 U74 ( .A(n244), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U75 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  XNOR2_X1 U76 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U77 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U78 ( .A(n240), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U79 ( .A1(n235), .A2(B[25]), .ZN(n240) );
  OR3_X1 U80 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U83 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U84 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U88 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U91 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U94 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U97 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U100 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U104 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U107 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR3_X1 U123 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_5 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_5_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_4_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n191, n192, n193, n194, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n190, n195, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U82 ( .A(n192), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U83 ( .A(n194), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n191), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n196), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n252), .ZN(n191) );
  OR3_X1 U2 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U5 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U6 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U7 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U8 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U9 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U10 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U11 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U12 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U13 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U14 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U15 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U16 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U17 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U19 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U20 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U21 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U22 ( .A(n209), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U23 ( .A1(n222), .A2(B[37]), .ZN(n209) );
  XNOR2_X1 U24 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U25 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U26 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U27 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U28 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U29 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U30 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U31 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U32 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U33 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  XNOR2_X1 U34 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U35 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U36 ( .A(n205), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U37 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  XNOR2_X1 U38 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U39 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  XNOR2_X1 U40 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U41 ( .A1(n191), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U42 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U43 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U44 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U45 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U46 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U47 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U48 ( .A(n215), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U49 ( .A1(n218), .A2(B[41]), .ZN(n215) );
  XNOR2_X1 U50 ( .A(n190), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U51 ( .A1(n214), .A2(B[45]), .ZN(n190) );
  XNOR2_X1 U52 ( .A(n195), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U53 ( .A1(n208), .A2(B[49]), .ZN(n195) );
  OR2_X1 U54 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  XNOR2_X1 U55 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U56 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U57 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U58 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U59 ( .A(B[8]), .B(n193), .ZN(DIFF[8]) );
  NOR2_X1 U60 ( .A1(B[7]), .A2(n194), .ZN(n193) );
  XNOR2_X1 U61 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U62 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U63 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U64 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U65 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U66 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U67 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U68 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U69 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U70 ( .A1(n196), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U71 ( .A(n227), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U72 ( .A1(n192), .A2(B[9]), .ZN(n227) );
  XNOR2_X1 U73 ( .A(n231), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U74 ( .A1(n247), .A2(B[13]), .ZN(n231) );
  XNOR2_X1 U75 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U76 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U77 ( .A(n236), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U78 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  XNOR2_X1 U79 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U80 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  OR3_X1 U81 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U84 ( .A1(B[10]), .A2(B[9]), .A3(n192), .ZN(n249) );
  OR3_X1 U91 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U94 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U97 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U100 ( .A1(B[5]), .A2(B[6]), .A3(n196), .ZN(n194) );
  OR3_X1 U104 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U107 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U110 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U113 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U116 ( .A1(B[7]), .A2(B[8]), .A3(n194), .ZN(n192) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n196) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_4 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_4_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_3_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U4 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  XNOR2_X1 U1 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U2 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U3 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U5 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U6 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U7 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  OR3_X1 U8 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  NAND2_X1 U9 ( .A1(n197), .A2(n252), .ZN(n196) );
  OR3_X1 U10 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  NOR3_X1 U11 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U12 ( .A(n223), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U13 ( .A1(n226), .A2(B[33]), .ZN(n223) );
  XNOR2_X1 U14 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U15 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U16 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U17 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U18 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U19 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U20 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U21 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U22 ( .A(n215), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U23 ( .A1(n204), .A2(B[53]), .ZN(n215) );
  XNOR2_X1 U24 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U25 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U26 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U27 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U28 ( .A(n209), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U29 ( .A1(n214), .A2(B[45]), .ZN(n209) );
  XNOR2_X1 U30 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U31 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U32 ( .A(n193), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U33 ( .A1(n200), .A2(B[57]), .ZN(n193) );
  XNOR2_X1 U34 ( .A(n205), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U35 ( .A1(n218), .A2(B[41]), .ZN(n205) );
  XNOR2_X1 U36 ( .A(n195), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U37 ( .A1(n222), .A2(B[37]), .ZN(n195) );
  OR3_X1 U38 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U39 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U40 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U41 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U42 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U43 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U44 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U45 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U46 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U47 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U48 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U49 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  NOR2_X1 U50 ( .A1(n230), .A2(B[29]), .ZN(n219) );
  XNOR2_X1 U51 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U52 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U53 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U54 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U55 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U56 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U57 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U58 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U61 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U62 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U63 ( .A(n227), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U64 ( .A1(n194), .A2(B[5]), .ZN(n227) );
  XNOR2_X1 U65 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U66 ( .A1(n190), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U67 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U68 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U69 ( .A(n248), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U70 ( .A1(n239), .A2(B[21]), .ZN(n248) );
  XNOR2_X1 U71 ( .A(n240), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U72 ( .A1(n235), .A2(B[25]), .ZN(n240) );
  XNOR2_X1 U73 ( .A(n244), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U74 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  XNOR2_X1 U75 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U76 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U77 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U78 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U79 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U80 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U83 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U84 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U88 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U91 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U94 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U97 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U100 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U104 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U107 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(n219), .B(B[30]), .ZN(DIFF[30]) );
  OR3_X1 U123 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_3 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_3_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_2_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n191, n192, n193, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n190, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n253;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U82 ( .A(n192), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U83 ( .A(n194), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n191), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n196), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n253), .ZN(n191) );
  OR3_X1 U2 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  OR3_X1 U4 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U7 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U8 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U9 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U10 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U11 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U12 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U13 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U14 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U15 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U16 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U17 ( .A(n223), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U18 ( .A1(n226), .A2(B[33]), .ZN(n223) );
  XNOR2_X1 U19 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U20 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U21 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U22 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U23 ( .A(n215), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U24 ( .A1(n218), .A2(B[41]), .ZN(n215) );
  XNOR2_X1 U25 ( .A(n190), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U26 ( .A1(n191), .A2(B[62]), .ZN(n190) );
  XNOR2_X1 U27 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U28 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U29 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U30 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U31 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U32 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U33 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U34 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U35 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U36 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U37 ( .A(n209), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U38 ( .A1(n214), .A2(B[45]), .ZN(n209) );
  XNOR2_X1 U39 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U40 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U41 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U42 ( .A(n205), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U43 ( .A1(n200), .A2(B[57]), .ZN(n205) );
  OR3_X1 U44 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U45 ( .A(n189), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U46 ( .A1(n230), .A2(B[29]), .ZN(n189) );
  XNOR2_X1 U47 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U48 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  XNOR2_X1 U49 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U50 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U51 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U52 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U53 ( .A(B[8]), .B(n193), .ZN(DIFF[8]) );
  NOR2_X1 U54 ( .A1(B[7]), .A2(n194), .ZN(n193) );
  XNOR2_X1 U55 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U56 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U57 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U58 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U59 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U60 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U61 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U62 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U63 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U64 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U65 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U66 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U67 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U68 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U69 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U70 ( .A1(n196), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U71 ( .A(n227), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U72 ( .A1(n192), .A2(B[9]), .ZN(n227) );
  XNOR2_X1 U73 ( .A(n231), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U74 ( .A1(n247), .A2(B[13]), .ZN(n231) );
  XNOR2_X1 U75 ( .A(n236), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U76 ( .A1(n243), .A2(B[17]), .ZN(n236) );
  XNOR2_X1 U77 ( .A(n240), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U78 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  XNOR2_X1 U79 ( .A(n244), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U80 ( .A1(n235), .A2(B[25]), .ZN(n244) );
  OR3_X1 U81 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U84 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U88 ( .A1(B[5]), .A2(B[6]), .A3(n196), .ZN(n194) );
  OR3_X1 U91 ( .A1(B[10]), .A2(B[9]), .A3(n192), .ZN(n249) );
  OR3_X1 U94 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U97 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U100 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U104 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U107 ( .A1(B[7]), .A2(B[8]), .A3(n194), .ZN(n192) );
  OR3_X1 U110 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U113 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U116 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n196) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n253) );
endmodule


module complement_NBIT64_2 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_2_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module complement_NBIT64_1_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n252;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U3 ( .A(n197), .B(n252), .Z(DIFF[61]) );
  XNOR2_X1 U1 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U2 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U4 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U5 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NAND2_X1 U6 ( .A1(n197), .A2(n252), .ZN(n196) );
  OR3_X1 U7 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U8 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U9 ( .A(n215), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U10 ( .A1(n226), .A2(B[33]), .ZN(n215) );
  NOR3_X1 U11 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U12 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U13 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U14 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U15 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U16 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U17 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U18 ( .A(n205), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U19 ( .A1(n208), .A2(B[49]), .ZN(n205) );
  XNOR2_X1 U20 ( .A(n193), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U21 ( .A1(n204), .A2(B[53]), .ZN(n193) );
  OR3_X1 U22 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U23 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U24 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U25 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U26 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U27 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U28 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U29 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U30 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U31 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U32 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U33 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U34 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U35 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U36 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U37 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U38 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U39 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U40 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U41 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U42 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  XNOR2_X1 U43 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U44 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U45 ( .A(n201), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U46 ( .A1(n214), .A2(B[45]), .ZN(n201) );
  NOR2_X1 U47 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U48 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U49 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U50 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U51 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U52 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U53 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U54 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U55 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U56 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U57 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U58 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U59 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U60 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U61 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U62 ( .A(n227), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U63 ( .A1(n194), .A2(B[5]), .ZN(n227) );
  XNOR2_X1 U64 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U65 ( .A1(n190), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U66 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U67 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U68 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U69 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  XNOR2_X1 U70 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U71 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U72 ( .A(n248), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U73 ( .A1(n235), .A2(B[25]), .ZN(n248) );
  XNOR2_X1 U74 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U75 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U76 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U77 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  OR3_X1 U78 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U79 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U80 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U83 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U84 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U88 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U91 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U94 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U97 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U100 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U104 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U107 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U110 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U113 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR3_X1 U123 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  INV_X1 U126 ( .A(B[61]), .ZN(n252) );
endmodule


module complement_NBIT64_1 ( A, Y );
  input [63:0] A;
  output [63:0] Y;


  complement_NBIT64_1_DW01_sub_0 sub_add_16_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module encoder_0 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n3, n4, n21, n18, n19, n20;

  AOI21_X2 U1 ( .B1(n19), .B2(n3), .A(n4), .ZN(Y[1]) );
  XOR2_X1 U7 ( .A(A[0]), .B(A[1]), .Z(n4) );
  AND2_X2 U2 ( .A1(n18), .A2(n4), .ZN(Y[0]) );
  AOI21_X1 U3 ( .B1(A[0]), .B2(A[1]), .A(n20), .ZN(Y[2]) );
  AOI21_X1 U4 ( .B1(A[0]), .B2(A[1]), .A(n20), .ZN(n21) );
  CLKBUF_X1 U5 ( .A(n20), .Z(n18) );
  NAND2_X1 U6 ( .A1(A[0]), .A2(n18), .ZN(n3) );
  INV_X1 U8 ( .A(A[2]), .ZN(n20) );
  INV_X1 U9 ( .A(n21), .ZN(n19) );
endmodule


module encoder_15 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n3, n4, n5, n18, n19;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n4) );
  AND2_X1 U1 ( .A1(n19), .A2(n4), .ZN(Y[0]) );
  NOR2_X1 U2 ( .A1(n19), .A2(n5), .ZN(Y[2]) );
  OR2_X1 U3 ( .A1(n19), .A2(n5), .ZN(n18) );
  AND2_X1 U4 ( .A1(A[1]), .A2(A[0]), .ZN(n5) );
  AOI21_X2 U5 ( .B1(n18), .B2(n3), .A(n4), .ZN(Y[1]) );
  NAND2_X1 U6 ( .A1(n5), .A2(n19), .ZN(n3) );
  INV_X1 U7 ( .A(A[2]), .ZN(n19) );
endmodule


module encoder_14 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n3, n4, n5, n16, n17;

  NOR2_X2 U3 ( .A1(n17), .A2(n5), .ZN(Y[2]) );
  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n4) );
  AOI21_X1 U1 ( .B1(n16), .B2(n3), .A(n4), .ZN(Y[1]) );
  NAND2_X1 U2 ( .A1(n5), .A2(n17), .ZN(n3) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n4), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n5) );
endmodule


module encoder_13 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n3, n4, n5, n16, n17;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n4) );
  NOR2_X1 U1 ( .A1(n17), .A2(n5), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n3), .A(n4), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n5), .A2(n17), .ZN(n3) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n4), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n5) );
endmodule


module encoder_12 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_11 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_10 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_9 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_8 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_7 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_6 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_5 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_4 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_3 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_2 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module encoder_1 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n16, n17, n19, n20, n21;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n20) );
  NOR2_X1 U1 ( .A1(n17), .A2(n19), .ZN(Y[2]) );
  AOI21_X1 U2 ( .B1(n16), .B2(n21), .A(n20), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n19), .A2(n17), .ZN(n21) );
  INV_X1 U4 ( .A(Y[2]), .ZN(n16) );
  AND2_X1 U5 ( .A1(n17), .A2(n20), .ZN(Y[0]) );
  INV_X1 U6 ( .A(A[2]), .ZN(n17) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n19) );
endmodule


module booth_encoder_NBIT32 ( A, Y );
  input [31:0] A;
  output [47:0] Y;


  encoder_0 ENCODER_N_0 ( .A({A[1:0], 1'b0}), .Y(Y[2:0]) );
  encoder_15 ENCODER_N_1 ( .A(A[3:1]), .Y(Y[5:3]) );
  encoder_14 ENCODER_N_2 ( .A(A[5:3]), .Y(Y[8:6]) );
  encoder_13 ENCODER_N_3 ( .A(A[7:5]), .Y(Y[11:9]) );
  encoder_12 ENCODER_N_4 ( .A(A[9:7]), .Y(Y[14:12]) );
  encoder_11 ENCODER_N_5 ( .A(A[11:9]), .Y(Y[17:15]) );
  encoder_10 ENCODER_N_6 ( .A(A[13:11]), .Y(Y[20:18]) );
  encoder_9 ENCODER_N_7 ( .A(A[15:13]), .Y(Y[23:21]) );
  encoder_8 ENCODER_N_8 ( .A(A[17:15]), .Y(Y[26:24]) );
  encoder_7 ENCODER_N_9 ( .A(A[19:17]), .Y(Y[29:27]) );
  encoder_6 ENCODER_N_10 ( .A(A[21:19]), .Y(Y[32:30]) );
  encoder_5 ENCODER_N_11 ( .A(A[23:21]), .Y(Y[35:33]) );
  encoder_4 ENCODER_N_12 ( .A(A[25:23]), .Y(Y[38:36]) );
  encoder_3 ENCODER_N_13 ( .A(A[27:25]), .Y(Y[41:39]) );
  encoder_2 ENCODER_N_14 ( .A(A[29:27]), .Y(Y[44:42]) );
  encoder_1 ENCODER_N_15 ( .A(A[31:29]), .Y(Y[47:45]) );
endmodule


module MUX81_GENERIC_NBIT64_0 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319;

  NOR3_X2 U322 ( .A1(n1318), .A2(SEL[0]), .A3(n1317), .ZN(n10) );
  NOR3_X2 U1 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1317), .ZN(n11) );
  BUF_X1 U2 ( .A(n14), .Z(n1269) );
  CLKBUF_X1 U3 ( .A(n10), .Z(n1303) );
  BUF_X1 U4 ( .A(n11), .Z(n1264) );
  BUF_X1 U5 ( .A(n8), .Z(n1265) );
  CLKBUF_X1 U6 ( .A(n10), .Z(n1301) );
  CLKBUF_X1 U7 ( .A(n1318), .Z(n1266) );
  CLKBUF_X3 U8 ( .A(n1269), .Z(n1280) );
  BUF_X1 U9 ( .A(n10), .Z(n1304) );
  CLKBUF_X3 U10 ( .A(n10), .Z(n1300) );
  CLKBUF_X3 U11 ( .A(n10), .Z(n1302) );
  CLKBUF_X3 U12 ( .A(n1269), .Z(n1279) );
  CLKBUF_X1 U13 ( .A(n1269), .Z(n1278) );
  CLKBUF_X3 U14 ( .A(n1265), .Z(n1315) );
  CLKBUF_X1 U15 ( .A(n8), .Z(n1313) );
  INV_X1 U16 ( .A(n1303), .ZN(n1267) );
  INV_X1 U17 ( .A(n1267), .ZN(n1268) );
  BUF_X2 U18 ( .A(n1264), .Z(n1295) );
  AOI22_X1 U19 ( .A1(G[37]), .A2(n1301), .B1(E[37]), .B2(n1296), .ZN(n150) );
  AOI22_X1 U20 ( .A1(G[32]), .A2(n1301), .B1(E[32]), .B2(n1296), .ZN(n170) );
  AOI22_X1 U21 ( .A1(G[36]), .A2(n1302), .B1(E[36]), .B2(n1296), .ZN(n154) );
  AOI22_X1 U22 ( .A1(G[40]), .A2(n1302), .B1(E[40]), .B2(n1296), .ZN(n134) );
  AOI22_X1 U23 ( .A1(G[41]), .A2(n1300), .B1(E[41]), .B2(n1296), .ZN(n130) );
  AOI22_X1 U24 ( .A1(G[54]), .A2(n1268), .B1(E[54]), .B2(n1298), .ZN(n74) );
  AOI22_X1 U25 ( .A1(G[39]), .A2(n1304), .B1(E[39]), .B2(n1296), .ZN(n142) );
  AOI22_X1 U26 ( .A1(G[55]), .A2(n1268), .B1(E[55]), .B2(n1298), .ZN(n70) );
  AOI22_X1 U27 ( .A1(G[56]), .A2(n1268), .B1(E[56]), .B2(n1298), .ZN(n66) );
  AOI22_X1 U28 ( .A1(G[57]), .A2(n1268), .B1(E[57]), .B2(n1298), .ZN(n62) );
  AOI22_X1 U29 ( .A1(G[60]), .A2(n1268), .B1(E[60]), .B2(n1298), .ZN(n50) );
  AOI22_X1 U30 ( .A1(G[58]), .A2(n1268), .B1(E[58]), .B2(n1298), .ZN(n58) );
  AOI22_X1 U31 ( .A1(G[63]), .A2(n1268), .B1(E[63]), .B2(n1298), .ZN(n38) );
  AOI22_X1 U32 ( .A1(G[61]), .A2(n1268), .B1(E[61]), .B2(n1298), .ZN(n46) );
  AOI22_X1 U33 ( .A1(G[62]), .A2(n1268), .B1(E[62]), .B2(n1298), .ZN(n42) );
  AOI22_X1 U34 ( .A1(G[59]), .A2(n1268), .B1(E[59]), .B2(n1298), .ZN(n54) );
  AOI22_X1 U35 ( .A1(G[42]), .A2(n1301), .B1(E[42]), .B2(n1296), .ZN(n126) );
  AOI22_X1 U36 ( .A1(G[34]), .A2(n1300), .B1(E[34]), .B2(n1296), .ZN(n162) );
  AOI22_X1 U37 ( .A1(G[38]), .A2(n1300), .B1(E[38]), .B2(n1296), .ZN(n146) );
  AOI22_X1 U38 ( .A1(G[35]), .A2(n1304), .B1(E[35]), .B2(n1296), .ZN(n158) );
  AOI22_X1 U39 ( .A1(G[33]), .A2(n1302), .B1(E[33]), .B2(n1296), .ZN(n166) );
  BUF_X1 U40 ( .A(n9), .Z(n1305) );
  BUF_X1 U41 ( .A(n9), .Z(n1306) );
  BUF_X1 U42 ( .A(n9), .Z(n1307) );
  BUF_X1 U43 ( .A(n9), .Z(n1308) );
  BUF_X1 U44 ( .A(n9), .Z(n1309) );
  CLKBUF_X1 U45 ( .A(n1265), .Z(n1311) );
  CLKBUF_X1 U46 ( .A(n1265), .Z(n1314) );
  CLKBUF_X1 U47 ( .A(n1265), .Z(n1312) );
  CLKBUF_X1 U48 ( .A(n1269), .Z(n1276) );
  BUF_X2 U49 ( .A(n11), .Z(n1296) );
  BUF_X2 U50 ( .A(n1264), .Z(n1294) );
  BUF_X2 U51 ( .A(n11), .Z(n1298) );
  AOI22_X1 U52 ( .A1(G[24]), .A2(n1302), .B1(E[24]), .B2(n1295), .ZN(n206) );
  AOI22_X1 U53 ( .A1(G[21]), .A2(n1302), .B1(E[21]), .B2(n1295), .ZN(n218) );
  AOI22_X1 U54 ( .A1(G[31]), .A2(n1300), .B1(E[31]), .B2(n1295), .ZN(n174) );
  AOI22_X1 U55 ( .A1(G[27]), .A2(n1302), .B1(E[27]), .B2(n1295), .ZN(n194) );
  AOI22_X1 U56 ( .A1(G[23]), .A2(n1304), .B1(E[23]), .B2(n1295), .ZN(n210) );
  AOI22_X1 U57 ( .A1(G[2]), .A2(n1302), .B1(E[2]), .B2(n1295), .ZN(n182) );
  AOI22_X1 U58 ( .A1(G[20]), .A2(n1300), .B1(E[20]), .B2(n1294), .ZN(n222) );
  AOI22_X1 U59 ( .A1(G[17]), .A2(n1302), .B1(E[17]), .B2(n1294), .ZN(n238) );
  AOI22_X1 U60 ( .A1(G[19]), .A2(n1301), .B1(E[19]), .B2(n1294), .ZN(n230) );
  AOI22_X1 U61 ( .A1(G[15]), .A2(n1302), .B1(E[15]), .B2(n1294), .ZN(n246) );
  AOI22_X1 U62 ( .A1(G[9]), .A2(n1301), .B1(E[9]), .B2(n1299), .ZN(n18) );
  BUF_X2 U63 ( .A(n11), .Z(n1297) );
  AOI22_X1 U64 ( .A1(G[13]), .A2(n1300), .B1(E[13]), .B2(n1294), .ZN(n254) );
  INV_X1 U65 ( .A(SEL[0]), .ZN(n1319) );
  BUF_X1 U66 ( .A(n12), .Z(n1289) );
  BUF_X1 U67 ( .A(n12), .Z(n1291) );
  BUF_X1 U68 ( .A(n12), .Z(n1288) );
  BUF_X1 U69 ( .A(n13), .Z(n1283) );
  BUF_X1 U70 ( .A(n13), .Z(n1285) );
  BUF_X1 U71 ( .A(n13), .Z(n1282) );
  BUF_X1 U72 ( .A(n15), .Z(n1270) );
  BUF_X1 U73 ( .A(n15), .Z(n1274) );
  BUF_X1 U74 ( .A(n12), .Z(n1290) );
  BUF_X1 U75 ( .A(n12), .Z(n1292) );
  BUF_X1 U76 ( .A(n15), .Z(n1271) );
  BUF_X1 U77 ( .A(n13), .Z(n1284) );
  BUF_X1 U78 ( .A(n13), .Z(n1286) );
  BUF_X1 U79 ( .A(n15), .Z(n1272) );
  BUF_X1 U80 ( .A(n15), .Z(n1273) );
  AOI22_X1 U81 ( .A1(G[14]), .A2(n1302), .B1(E[14]), .B2(n1294), .ZN(n250) );
  AOI22_X1 U82 ( .A1(G[28]), .A2(n1304), .B1(E[28]), .B2(n1295), .ZN(n190) );
  AOI22_X1 U83 ( .A1(G[26]), .A2(n1300), .B1(E[26]), .B2(n1295), .ZN(n198) );
  AOI22_X1 U84 ( .A1(G[30]), .A2(n1302), .B1(E[30]), .B2(n1295), .ZN(n178) );
  AOI22_X1 U85 ( .A1(G[22]), .A2(n1301), .B1(E[22]), .B2(n1295), .ZN(n214) );
  AOI22_X1 U86 ( .A1(G[18]), .A2(n1304), .B1(E[18]), .B2(n1294), .ZN(n234) );
  AOI22_X1 U87 ( .A1(G[16]), .A2(n1300), .B1(E[16]), .B2(n1294), .ZN(n242) );
  AOI22_X1 U88 ( .A1(G[12]), .A2(n1300), .B1(E[12]), .B2(n1294), .ZN(n258) );
  AOI22_X1 U89 ( .A1(G[8]), .A2(n1300), .B1(E[8]), .B2(n1299), .ZN(n26) );
  AOI22_X1 U90 ( .A1(G[25]), .A2(n1301), .B1(E[25]), .B2(n1295), .ZN(n202) );
  AOI22_X1 U91 ( .A1(G[29]), .A2(n1300), .B1(E[29]), .B2(n1295), .ZN(n186) );
  AOI22_X1 U92 ( .A1(C[7]), .A2(n1277), .B1(A[7]), .B2(n1274), .ZN(n28) );
  AOI22_X1 U93 ( .A1(F[4]), .A2(n1291), .B1(D[4]), .B2(n1285), .ZN(n93) );
  NAND4_X1 U94 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(Y[8]) );
  AOI22_X1 U95 ( .A1(F[8]), .A2(n1293), .B1(D[8]), .B2(n1287), .ZN(n25) );
  AOI22_X1 U96 ( .A1(B[8]), .A2(n1315), .B1(H[8]), .B2(n1310), .ZN(n27) );
  AOI22_X1 U97 ( .A1(C[8]), .A2(n1280), .B1(A[8]), .B2(n1275), .ZN(n24) );
  NAND4_X1 U98 ( .A1(n180), .A2(n181), .A3(n182), .A4(n183), .ZN(Y[2]) );
  AOI22_X1 U99 ( .A1(F[2]), .A2(n1289), .B1(D[2]), .B2(n1283), .ZN(n181) );
  AOI22_X1 U100 ( .A1(B[2]), .A2(n1313), .B1(H[2]), .B2(n1306), .ZN(n183) );
  AOI22_X1 U101 ( .A1(F[38]), .A2(n1290), .B1(D[38]), .B2(n1284), .ZN(n145) );
  AOI22_X1 U102 ( .A1(B[38]), .A2(n1315), .B1(H[38]), .B2(n1307), .ZN(n147) );
  AOI22_X1 U103 ( .A1(F[11]), .A2(n1288), .B1(D[11]), .B2(n1282), .ZN(n261) );
  AOI22_X1 U104 ( .A1(B[11]), .A2(n1316), .B1(H[11]), .B2(n1305), .ZN(n263) );
  AOI22_X1 U105 ( .A1(C[11]), .A2(n1280), .B1(A[11]), .B2(n1270), .ZN(n260) );
  AOI22_X1 U106 ( .A1(F[5]), .A2(n1293), .B1(D[5]), .B2(n1287), .ZN(n21) );
  AOI22_X1 U107 ( .A1(B[5]), .A2(n1313), .B1(H[5]), .B2(n1310), .ZN(n23) );
  AOI22_X1 U108 ( .A1(F[10]), .A2(n1293), .B1(D[10]), .B2(n1287), .ZN(n5) );
  AOI22_X1 U109 ( .A1(B[10]), .A2(n1314), .B1(H[10]), .B2(n1310), .ZN(n7) );
  AOI22_X1 U110 ( .A1(C[10]), .A2(n1277), .B1(A[10]), .B2(n1275), .ZN(n4) );
  AOI22_X1 U111 ( .A1(F[35]), .A2(n1290), .B1(D[35]), .B2(n1284), .ZN(n157) );
  AOI22_X1 U112 ( .A1(B[35]), .A2(n1314), .B1(H[35]), .B2(n1307), .ZN(n159) );
  AOI22_X1 U113 ( .A1(F[43]), .A2(n1291), .B1(D[43]), .B2(n1285), .ZN(n121) );
  AOI22_X1 U114 ( .A1(B[43]), .A2(n1312), .B1(H[43]), .B2(n1308), .ZN(n123) );
  NAND4_X1 U115 ( .A1(n252), .A2(n253), .A3(n254), .A4(n255), .ZN(Y[13]) );
  AOI22_X1 U116 ( .A1(F[13]), .A2(n1288), .B1(D[13]), .B2(n1282), .ZN(n253) );
  AOI22_X1 U117 ( .A1(B[13]), .A2(n1311), .B1(H[13]), .B2(n1305), .ZN(n255) );
  AOI22_X1 U118 ( .A1(C[13]), .A2(n1277), .B1(A[13]), .B2(n1270), .ZN(n252) );
  AOI22_X1 U119 ( .A1(C[6]), .A2(n1278), .B1(A[6]), .B2(n1274), .ZN(n32) );
  NAND4_X1 U120 ( .A1(n244), .A2(n245), .A3(n246), .A4(n247), .ZN(Y[15]) );
  AOI22_X1 U121 ( .A1(F[15]), .A2(n1288), .B1(D[15]), .B2(n1282), .ZN(n245) );
  AOI22_X1 U122 ( .A1(B[15]), .A2(n1316), .B1(H[15]), .B2(n1305), .ZN(n247) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n1280), .B1(A[15]), .B2(n1270), .ZN(n244) );
  NAND4_X1 U124 ( .A1(n164), .A2(n165), .A3(n166), .A4(n167), .ZN(Y[33]) );
  AOI22_X1 U125 ( .A1(F[33]), .A2(n1290), .B1(D[33]), .B2(n1284), .ZN(n165) );
  AOI22_X1 U126 ( .A1(B[33]), .A2(n1311), .B1(H[33]), .B2(n1307), .ZN(n167) );
  NAND4_X1 U127 ( .A1(n168), .A2(n169), .A3(n170), .A4(n171), .ZN(Y[32]) );
  AOI22_X1 U128 ( .A1(F[32]), .A2(n1290), .B1(D[32]), .B2(n1284), .ZN(n169) );
  AOI22_X1 U129 ( .A1(B[32]), .A2(n1312), .B1(H[32]), .B2(n1307), .ZN(n171) );
  NAND4_X1 U130 ( .A1(n148), .A2(n149), .A3(n150), .A4(n151), .ZN(Y[37]) );
  AOI22_X1 U131 ( .A1(F[37]), .A2(n1290), .B1(D[37]), .B2(n1284), .ZN(n149) );
  AOI22_X1 U132 ( .A1(B[37]), .A2(n1312), .B1(H[37]), .B2(n1307), .ZN(n151) );
  NAND4_X1 U133 ( .A1(n152), .A2(n153), .A3(n154), .A4(n155), .ZN(Y[36]) );
  AOI22_X1 U134 ( .A1(F[36]), .A2(n1290), .B1(D[36]), .B2(n1284), .ZN(n153) );
  AOI22_X1 U135 ( .A1(B[36]), .A2(n1315), .B1(H[36]), .B2(n1307), .ZN(n155) );
  NAND4_X1 U136 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(Y[34]) );
  AOI22_X1 U137 ( .A1(F[34]), .A2(n1290), .B1(D[34]), .B2(n1284), .ZN(n161) );
  AOI22_X1 U138 ( .A1(B[34]), .A2(n1316), .B1(H[34]), .B2(n1307), .ZN(n163) );
  NAND4_X1 U139 ( .A1(n132), .A2(n133), .A3(n134), .A4(n135), .ZN(Y[40]) );
  AOI22_X1 U140 ( .A1(F[40]), .A2(n1290), .B1(D[40]), .B2(n1284), .ZN(n133) );
  AOI22_X1 U141 ( .A1(B[40]), .A2(n1316), .B1(H[40]), .B2(n1307), .ZN(n135) );
  NAND4_X1 U142 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(Y[52]) );
  AOI22_X1 U143 ( .A1(F[52]), .A2(n1291), .B1(D[52]), .B2(n1285), .ZN(n81) );
  AOI22_X1 U144 ( .A1(B[52]), .A2(n1315), .B1(H[52]), .B2(n1308), .ZN(n83) );
  NAND4_X1 U145 ( .A1(n100), .A2(n101), .A3(n102), .A4(n103), .ZN(Y[48]) );
  AOI22_X1 U146 ( .A1(F[48]), .A2(n1291), .B1(D[48]), .B2(n1285), .ZN(n101) );
  AOI22_X1 U147 ( .A1(B[48]), .A2(n1312), .B1(H[48]), .B2(n1308), .ZN(n103) );
  NAND4_X1 U148 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(Y[53]) );
  AOI22_X1 U149 ( .A1(F[53]), .A2(n1291), .B1(D[53]), .B2(n1285), .ZN(n77) );
  AOI22_X1 U150 ( .A1(B[53]), .A2(n1315), .B1(H[53]), .B2(n1308), .ZN(n79) );
  NAND4_X1 U151 ( .A1(n96), .A2(n97), .A3(n98), .A4(n99), .ZN(Y[49]) );
  AOI22_X1 U152 ( .A1(F[49]), .A2(n1291), .B1(D[49]), .B2(n1285), .ZN(n97) );
  AOI22_X1 U153 ( .A1(B[49]), .A2(n1311), .B1(H[49]), .B2(n1308), .ZN(n99) );
  NAND4_X1 U154 ( .A1(n88), .A2(n89), .A3(n90), .A4(n91), .ZN(Y[50]) );
  AOI22_X1 U155 ( .A1(F[50]), .A2(n1291), .B1(D[50]), .B2(n1285), .ZN(n89) );
  AOI22_X1 U156 ( .A1(B[50]), .A2(n1316), .B1(H[50]), .B2(n1308), .ZN(n91) );
  NAND4_X1 U157 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(Y[41]) );
  AOI22_X1 U158 ( .A1(F[41]), .A2(n1290), .B1(D[41]), .B2(n1284), .ZN(n129) );
  AOI22_X1 U159 ( .A1(B[41]), .A2(n1314), .B1(H[41]), .B2(n1307), .ZN(n131) );
  NAND4_X1 U160 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(Y[44]) );
  AOI22_X1 U161 ( .A1(F[44]), .A2(n1291), .B1(D[44]), .B2(n1285), .ZN(n117) );
  AOI22_X1 U162 ( .A1(B[44]), .A2(n1311), .B1(H[44]), .B2(n1308), .ZN(n119) );
  NAND4_X1 U163 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(Y[45]) );
  AOI22_X1 U164 ( .A1(F[45]), .A2(n1291), .B1(D[45]), .B2(n1285), .ZN(n113) );
  AOI22_X1 U165 ( .A1(B[45]), .A2(n1316), .B1(H[45]), .B2(n1308), .ZN(n115) );
  NAND4_X1 U166 ( .A1(n124), .A2(n125), .A3(n126), .A4(n127), .ZN(Y[42]) );
  AOI22_X1 U167 ( .A1(F[42]), .A2(n1290), .B1(D[42]), .B2(n1284), .ZN(n125) );
  AOI22_X1 U168 ( .A1(B[42]), .A2(n1315), .B1(H[42]), .B2(n1307), .ZN(n127) );
  NAND4_X1 U169 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(Y[46]) );
  AOI22_X1 U170 ( .A1(F[46]), .A2(n1291), .B1(D[46]), .B2(n1285), .ZN(n109) );
  AOI22_X1 U171 ( .A1(B[46]), .A2(n1314), .B1(H[46]), .B2(n1308), .ZN(n111) );
  NAND4_X1 U172 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(Y[47]) );
  AOI22_X1 U173 ( .A1(F[47]), .A2(n1291), .B1(D[47]), .B2(n1285), .ZN(n105) );
  AOI22_X1 U174 ( .A1(B[47]), .A2(n1315), .B1(H[47]), .B2(n1308), .ZN(n107) );
  AOI22_X1 U175 ( .A1(B[4]), .A2(n1313), .B1(H[4]), .B2(n1308), .ZN(n95) );
  AOI22_X1 U176 ( .A1(B[3]), .A2(n1313), .B1(H[3]), .B2(n1307), .ZN(n139) );
  NAND4_X1 U177 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(Y[6]) );
  AOI22_X1 U178 ( .A1(F[6]), .A2(n1292), .B1(D[6]), .B2(n1286), .ZN(n33) );
  AOI22_X1 U179 ( .A1(B[6]), .A2(n1313), .B1(H[6]), .B2(n1309), .ZN(n35) );
  AOI22_X1 U180 ( .A1(G[6]), .A2(n1303), .B1(E[6]), .B2(n1298), .ZN(n34) );
  NAND4_X1 U181 ( .A1(n220), .A2(n221), .A3(n222), .A4(n223), .ZN(Y[20]) );
  AOI22_X1 U182 ( .A1(F[20]), .A2(n1288), .B1(D[20]), .B2(n1282), .ZN(n221) );
  AOI22_X1 U183 ( .A1(B[20]), .A2(n1314), .B1(H[20]), .B2(n1305), .ZN(n223) );
  AOI22_X1 U184 ( .A1(C[20]), .A2(n1279), .B1(A[20]), .B2(n1270), .ZN(n220) );
  NAND4_X1 U185 ( .A1(n232), .A2(n233), .A3(n234), .A4(n235), .ZN(Y[18]) );
  AOI22_X1 U186 ( .A1(F[18]), .A2(n1288), .B1(D[18]), .B2(n1282), .ZN(n233) );
  AOI22_X1 U187 ( .A1(B[18]), .A2(n1311), .B1(H[18]), .B2(n1305), .ZN(n235) );
  AOI22_X1 U188 ( .A1(C[18]), .A2(n1277), .B1(A[18]), .B2(n1270), .ZN(n232) );
  NAND4_X1 U189 ( .A1(n228), .A2(n229), .A3(n230), .A4(n231), .ZN(Y[19]) );
  AOI22_X1 U190 ( .A1(F[19]), .A2(n1288), .B1(D[19]), .B2(n1282), .ZN(n229) );
  AOI22_X1 U191 ( .A1(B[19]), .A2(n1316), .B1(H[19]), .B2(n1305), .ZN(n231) );
  AOI22_X1 U192 ( .A1(C[19]), .A2(n1280), .B1(A[19]), .B2(n1270), .ZN(n228) );
  NAND4_X1 U193 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(Y[12]) );
  AOI22_X1 U194 ( .A1(F[12]), .A2(n1288), .B1(D[12]), .B2(n1282), .ZN(n257) );
  AOI22_X1 U195 ( .A1(B[12]), .A2(n1314), .B1(H[12]), .B2(n1305), .ZN(n259) );
  AOI22_X1 U196 ( .A1(C[12]), .A2(n1279), .B1(A[12]), .B2(n1270), .ZN(n256) );
  NAND4_X1 U197 ( .A1(n248), .A2(n249), .A3(n250), .A4(n251), .ZN(Y[14]) );
  AOI22_X1 U198 ( .A1(F[14]), .A2(n1288), .B1(D[14]), .B2(n1282), .ZN(n249) );
  AOI22_X1 U199 ( .A1(B[14]), .A2(n1312), .B1(H[14]), .B2(n1305), .ZN(n251) );
  AOI22_X1 U200 ( .A1(C[14]), .A2(n1279), .B1(A[14]), .B2(n1270), .ZN(n248) );
  NAND4_X1 U201 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(Y[54]) );
  AOI22_X1 U202 ( .A1(F[54]), .A2(n1292), .B1(D[54]), .B2(n1286), .ZN(n73) );
  AOI22_X1 U203 ( .A1(B[54]), .A2(n1311), .B1(H[54]), .B2(n1309), .ZN(n75) );
  AOI22_X1 U204 ( .A1(C[54]), .A2(n1280), .B1(A[54]), .B2(n1274), .ZN(n72) );
  NAND4_X1 U205 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(Y[56]) );
  AOI22_X1 U206 ( .A1(F[56]), .A2(n1292), .B1(D[56]), .B2(n1286), .ZN(n65) );
  AOI22_X1 U207 ( .A1(B[56]), .A2(n1316), .B1(H[56]), .B2(n1309), .ZN(n67) );
  AOI22_X1 U208 ( .A1(C[56]), .A2(n1277), .B1(A[56]), .B2(n1274), .ZN(n64) );
  NAND4_X1 U209 ( .A1(n60), .A2(n61), .A3(n62), .A4(n63), .ZN(Y[57]) );
  AOI22_X1 U210 ( .A1(F[57]), .A2(n1292), .B1(D[57]), .B2(n1286), .ZN(n61) );
  AOI22_X1 U211 ( .A1(B[57]), .A2(n1314), .B1(H[57]), .B2(n1309), .ZN(n63) );
  AOI22_X1 U212 ( .A1(C[57]), .A2(n1280), .B1(A[57]), .B2(n1274), .ZN(n60) );
  NAND4_X1 U213 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .ZN(Y[60]) );
  AOI22_X1 U214 ( .A1(F[60]), .A2(n1292), .B1(D[60]), .B2(n1286), .ZN(n49) );
  AOI22_X1 U215 ( .A1(B[60]), .A2(n1311), .B1(H[60]), .B2(n1309), .ZN(n51) );
  AOI22_X1 U216 ( .A1(C[60]), .A2(n1281), .B1(A[60]), .B2(n1274), .ZN(n48) );
  NAND4_X1 U217 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(Y[58]) );
  AOI22_X1 U218 ( .A1(F[58]), .A2(n1292), .B1(D[58]), .B2(n1286), .ZN(n57) );
  AOI22_X1 U219 ( .A1(B[58]), .A2(n1312), .B1(H[58]), .B2(n1309), .ZN(n59) );
  AOI22_X1 U220 ( .A1(C[58]), .A2(n1276), .B1(A[58]), .B2(n1274), .ZN(n56) );
  NAND4_X1 U221 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(Y[61]) );
  AOI22_X1 U222 ( .A1(F[61]), .A2(n1292), .B1(D[61]), .B2(n1286), .ZN(n45) );
  AOI22_X1 U223 ( .A1(B[61]), .A2(n1315), .B1(H[61]), .B2(n1309), .ZN(n47) );
  AOI22_X1 U224 ( .A1(C[61]), .A2(n1277), .B1(A[61]), .B2(n1274), .ZN(n44) );
  NAND4_X1 U225 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(Y[62]) );
  AOI22_X1 U226 ( .A1(F[62]), .A2(n1292), .B1(D[62]), .B2(n1286), .ZN(n41) );
  AOI22_X1 U227 ( .A1(B[62]), .A2(n1315), .B1(H[62]), .B2(n1309), .ZN(n43) );
  AOI22_X1 U228 ( .A1(C[62]), .A2(n1280), .B1(A[62]), .B2(n1274), .ZN(n40) );
  NAND4_X1 U229 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(Y[63]) );
  AOI22_X1 U230 ( .A1(F[63]), .A2(n1292), .B1(D[63]), .B2(n1286), .ZN(n37) );
  AOI22_X1 U231 ( .A1(B[63]), .A2(n1315), .B1(H[63]), .B2(n1309), .ZN(n39) );
  AOI22_X1 U232 ( .A1(C[63]), .A2(n1276), .B1(A[63]), .B2(n1274), .ZN(n36) );
  NAND4_X1 U233 ( .A1(n216), .A2(n217), .A3(n218), .A4(n219), .ZN(Y[21]) );
  AOI22_X1 U234 ( .A1(F[21]), .A2(n1289), .B1(D[21]), .B2(n1283), .ZN(n217) );
  AOI22_X1 U235 ( .A1(B[21]), .A2(n1315), .B1(H[21]), .B2(n1306), .ZN(n219) );
  AOI22_X1 U236 ( .A1(C[21]), .A2(n1280), .B1(A[21]), .B2(n1271), .ZN(n216) );
  NAND4_X1 U237 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(Y[28]) );
  AOI22_X1 U238 ( .A1(F[28]), .A2(n1289), .B1(D[28]), .B2(n1283), .ZN(n189) );
  AOI22_X1 U239 ( .A1(B[28]), .A2(n1315), .B1(H[28]), .B2(n1306), .ZN(n191) );
  AOI22_X1 U240 ( .A1(C[28]), .A2(n1279), .B1(A[28]), .B2(n1271), .ZN(n188) );
  NAND4_X1 U241 ( .A1(n204), .A2(n205), .A3(n206), .A4(n207), .ZN(Y[24]) );
  AOI22_X1 U242 ( .A1(F[24]), .A2(n1289), .B1(D[24]), .B2(n1283), .ZN(n205) );
  AOI22_X1 U243 ( .A1(B[24]), .A2(n1315), .B1(H[24]), .B2(n1306), .ZN(n207) );
  AOI22_X1 U244 ( .A1(C[24]), .A2(n1277), .B1(A[24]), .B2(n1271), .ZN(n204) );
  NAND4_X1 U245 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(Y[25]) );
  AOI22_X1 U246 ( .A1(F[25]), .A2(n1289), .B1(D[25]), .B2(n1283), .ZN(n201) );
  AOI22_X1 U247 ( .A1(B[25]), .A2(n1311), .B1(H[25]), .B2(n1306), .ZN(n203) );
  AOI22_X1 U248 ( .A1(C[25]), .A2(n1279), .B1(A[25]), .B2(n1271), .ZN(n200) );
  NAND4_X1 U249 ( .A1(n212), .A2(n213), .A3(n214), .A4(n215), .ZN(Y[22]) );
  AOI22_X1 U250 ( .A1(F[22]), .A2(n1289), .B1(D[22]), .B2(n1283), .ZN(n213) );
  AOI22_X1 U251 ( .A1(B[22]), .A2(n1315), .B1(H[22]), .B2(n1306), .ZN(n215) );
  AOI22_X1 U252 ( .A1(C[22]), .A2(n1277), .B1(A[22]), .B2(n1271), .ZN(n212) );
  NAND4_X1 U253 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(Y[30]) );
  AOI22_X1 U254 ( .A1(F[30]), .A2(n1289), .B1(D[30]), .B2(n1283), .ZN(n177) );
  AOI22_X1 U255 ( .A1(B[30]), .A2(n1315), .B1(H[30]), .B2(n1306), .ZN(n179) );
  AOI22_X1 U256 ( .A1(C[30]), .A2(n1277), .B1(A[30]), .B2(n1271), .ZN(n176) );
  NAND4_X1 U257 ( .A1(n208), .A2(n209), .A3(n210), .A4(n211), .ZN(Y[23]) );
  AOI22_X1 U258 ( .A1(F[23]), .A2(n1289), .B1(D[23]), .B2(n1283), .ZN(n209) );
  AOI22_X1 U259 ( .A1(B[23]), .A2(n1312), .B1(H[23]), .B2(n1306), .ZN(n211) );
  AOI22_X1 U260 ( .A1(C[23]), .A2(n1279), .B1(A[23]), .B2(n1271), .ZN(n208) );
  NAND4_X1 U261 ( .A1(n19), .A2(n17), .A3(n18), .A4(n16), .ZN(Y[9]) );
  AOI22_X1 U262 ( .A1(F[9]), .A2(n1293), .B1(D[9]), .B2(n1287), .ZN(n17) );
  AOI22_X1 U263 ( .A1(B[9]), .A2(n1315), .B1(H[9]), .B2(n1310), .ZN(n19) );
  AOI22_X1 U264 ( .A1(C[9]), .A2(n1279), .B1(A[9]), .B2(n1275), .ZN(n16) );
  AOI22_X1 U265 ( .A1(C[5]), .A2(n1278), .B1(A[5]), .B2(n1275), .ZN(n20) );
  NAND4_X1 U266 ( .A1(n84), .A2(n85), .A3(n86), .A4(n87), .ZN(Y[51]) );
  AOI22_X1 U267 ( .A1(F[51]), .A2(n1291), .B1(D[51]), .B2(n1285), .ZN(n85) );
  AOI22_X1 U268 ( .A1(B[51]), .A2(n1314), .B1(H[51]), .B2(n1308), .ZN(n87) );
  NAND4_X1 U269 ( .A1(n68), .A2(n69), .A3(n70), .A4(n71), .ZN(Y[55]) );
  AOI22_X1 U270 ( .A1(F[55]), .A2(n1292), .B1(D[55]), .B2(n1286), .ZN(n69) );
  AOI22_X1 U271 ( .A1(B[55]), .A2(n1312), .B1(H[55]), .B2(n1309), .ZN(n71) );
  AOI22_X1 U272 ( .A1(C[55]), .A2(n1279), .B1(A[55]), .B2(n1274), .ZN(n68) );
  NAND4_X1 U273 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(Y[59]) );
  AOI22_X1 U274 ( .A1(F[59]), .A2(n1292), .B1(D[59]), .B2(n1286), .ZN(n53) );
  AOI22_X1 U275 ( .A1(B[59]), .A2(n1315), .B1(H[59]), .B2(n1309), .ZN(n55) );
  AOI22_X1 U276 ( .A1(C[59]), .A2(n1279), .B1(A[59]), .B2(n1274), .ZN(n52) );
  NAND4_X1 U277 ( .A1(n240), .A2(n241), .A3(n242), .A4(n243), .ZN(Y[16]) );
  AOI22_X1 U278 ( .A1(F[16]), .A2(n1288), .B1(D[16]), .B2(n1282), .ZN(n241) );
  AOI22_X1 U279 ( .A1(B[16]), .A2(n1315), .B1(H[16]), .B2(n1305), .ZN(n243) );
  AOI22_X1 U280 ( .A1(C[16]), .A2(n1276), .B1(A[16]), .B2(n1270), .ZN(n240) );
  NAND4_X1 U281 ( .A1(n238), .A2(n237), .A3(n236), .A4(n239), .ZN(Y[17]) );
  AOI22_X1 U282 ( .A1(F[17]), .A2(n1288), .B1(D[17]), .B2(n1282), .ZN(n237) );
  AOI22_X1 U283 ( .A1(B[17]), .A2(n1312), .B1(H[17]), .B2(n1305), .ZN(n239) );
  AOI22_X1 U284 ( .A1(C[17]), .A2(n1281), .B1(A[17]), .B2(n1270), .ZN(n236) );
  NAND4_X1 U285 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(Y[31]) );
  AOI22_X1 U286 ( .A1(F[31]), .A2(n1289), .B1(D[31]), .B2(n1283), .ZN(n173) );
  AOI22_X1 U287 ( .A1(B[31]), .A2(n1315), .B1(H[31]), .B2(n1306), .ZN(n175) );
  AOI22_X1 U288 ( .A1(C[31]), .A2(n1280), .B1(A[31]), .B2(n1271), .ZN(n172) );
  NAND4_X1 U289 ( .A1(n192), .A2(n193), .A3(n194), .A4(n195), .ZN(Y[27]) );
  AOI22_X1 U290 ( .A1(F[27]), .A2(n1289), .B1(D[27]), .B2(n1283), .ZN(n193) );
  AOI22_X1 U291 ( .A1(B[27]), .A2(n1316), .B1(H[27]), .B2(n1306), .ZN(n195) );
  AOI22_X1 U292 ( .A1(C[27]), .A2(n1277), .B1(A[27]), .B2(n1271), .ZN(n192) );
  NAND4_X1 U293 ( .A1(n140), .A2(n141), .A3(n142), .A4(n143), .ZN(Y[39]) );
  AOI22_X1 U294 ( .A1(F[39]), .A2(n1290), .B1(D[39]), .B2(n1284), .ZN(n141) );
  AOI22_X1 U295 ( .A1(B[39]), .A2(n1311), .B1(H[39]), .B2(n1307), .ZN(n143) );
  NAND4_X1 U296 ( .A1(n186), .A2(n185), .A3(n184), .A4(n187), .ZN(Y[29]) );
  AOI22_X1 U297 ( .A1(F[29]), .A2(n1289), .B1(D[29]), .B2(n1283), .ZN(n185) );
  AOI22_X1 U298 ( .A1(B[29]), .A2(n1314), .B1(H[29]), .B2(n1306), .ZN(n187) );
  AOI22_X1 U299 ( .A1(C[29]), .A2(n1280), .B1(A[29]), .B2(n1271), .ZN(n184) );
  NAND4_X1 U300 ( .A1(n196), .A2(n197), .A3(n198), .A4(n199), .ZN(Y[26]) );
  AOI22_X1 U301 ( .A1(F[26]), .A2(n1289), .B1(D[26]), .B2(n1283), .ZN(n197) );
  AOI22_X1 U302 ( .A1(B[26]), .A2(n1315), .B1(H[26]), .B2(n1306), .ZN(n199) );
  AOI22_X1 U303 ( .A1(C[26]), .A2(n1280), .B1(A[26]), .B2(n1271), .ZN(n196) );
  AOI22_X1 U304 ( .A1(C[1]), .A2(n1281), .B1(A[1]), .B2(n1270), .ZN(n224) );
  NAND4_X1 U305 ( .A1(n224), .A2(n225), .A3(n226), .A4(n227), .ZN(Y[1]) );
  AOI22_X1 U306 ( .A1(F[1]), .A2(n1288), .B1(D[1]), .B2(n1282), .ZN(n225) );
  AOI22_X1 U307 ( .A1(B[1]), .A2(n1316), .B1(H[1]), .B2(n1305), .ZN(n227) );
  AOI22_X1 U308 ( .A1(G[1]), .A2(n1304), .B1(E[1]), .B2(n1294), .ZN(n226) );
  AOI22_X1 U309 ( .A1(B[0]), .A2(n1314), .B1(H[0]), .B2(n1305), .ZN(n267) );
  NAND4_X1 U310 ( .A1(n264), .A2(n265), .A3(n266), .A4(n267), .ZN(Y[0]) );
  AOI22_X1 U311 ( .A1(C[0]), .A2(n1279), .B1(A[0]), .B2(n1270), .ZN(n264) );
  AOI22_X1 U312 ( .A1(F[0]), .A2(n1288), .B1(D[0]), .B2(n1282), .ZN(n265) );
  AOI22_X1 U313 ( .A1(G[0]), .A2(n1304), .B1(E[0]), .B2(n1294), .ZN(n266) );
  NAND4_X1 U314 ( .A1(n158), .A2(n157), .A3(n156), .A4(n159), .ZN(Y[35]) );
  NOR3_X1 U315 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1318), .ZN(n14) );
  AOI22_X1 U316 ( .A1(G[5]), .A2(n1300), .B1(E[5]), .B2(n1299), .ZN(n22) );
  AOI22_X1 U317 ( .A1(B[7]), .A2(n1313), .B1(H[7]), .B2(n1309), .ZN(n31) );
  NAND4_X1 U318 ( .A1(n22), .A2(n21), .A3(n20), .A4(n23), .ZN(Y[5]) );
  NAND4_X1 U319 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(Y[10]) );
  AOI22_X1 U320 ( .A1(F[3]), .A2(n1290), .B1(D[3]), .B2(n1284), .ZN(n137) );
  AOI22_X1 U321 ( .A1(G[3]), .A2(n1304), .B1(E[3]), .B2(n1296), .ZN(n138) );
  NOR3_X1 U323 ( .A1(n1266), .A2(n1319), .A3(n1317), .ZN(n9) );
  NAND4_X1 U324 ( .A1(n120), .A2(n121), .A3(n122), .A4(n123), .ZN(Y[43]) );
  AOI22_X1 U325 ( .A1(G[53]), .A2(n1268), .B1(E[53]), .B2(n1297), .ZN(n78) );
  AOI22_X1 U326 ( .A1(G[52]), .A2(n1268), .B1(E[52]), .B2(n1297), .ZN(n82) );
  AOI22_X1 U327 ( .A1(G[51]), .A2(n1268), .B1(E[51]), .B2(n1297), .ZN(n86) );
  AOI22_X1 U328 ( .A1(G[50]), .A2(n1268), .B1(E[50]), .B2(n1297), .ZN(n90) );
  AOI22_X1 U329 ( .A1(G[49]), .A2(n1268), .B1(E[49]), .B2(n1297), .ZN(n98) );
  AOI22_X1 U330 ( .A1(G[48]), .A2(n1268), .B1(E[48]), .B2(n1297), .ZN(n102) );
  AOI22_X1 U331 ( .A1(G[47]), .A2(n1268), .B1(E[47]), .B2(n1297), .ZN(n106) );
  AOI22_X1 U332 ( .A1(G[46]), .A2(n1268), .B1(E[46]), .B2(n1297), .ZN(n110) );
  AOI22_X1 U333 ( .A1(G[45]), .A2(n1268), .B1(E[45]), .B2(n1297), .ZN(n114) );
  AOI22_X1 U334 ( .A1(G[44]), .A2(n1268), .B1(E[44]), .B2(n1297), .ZN(n118) );
  AOI22_X1 U335 ( .A1(G[43]), .A2(n1268), .B1(E[43]), .B2(n1297), .ZN(n122) );
  NAND4_X1 U336 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(Y[4]) );
  AOI22_X1 U337 ( .A1(G[4]), .A2(n1303), .B1(E[4]), .B2(n1297), .ZN(n94) );
  AOI22_X1 U338 ( .A1(C[53]), .A2(n1277), .B1(A[53]), .B2(n1273), .ZN(n76) );
  AOI22_X1 U339 ( .A1(C[52]), .A2(n1281), .B1(A[52]), .B2(n1273), .ZN(n80) );
  AOI22_X1 U340 ( .A1(C[51]), .A2(n1276), .B1(A[51]), .B2(n1273), .ZN(n84) );
  AOI22_X1 U341 ( .A1(C[50]), .A2(n1279), .B1(A[50]), .B2(n1273), .ZN(n88) );
  AOI22_X1 U342 ( .A1(C[49]), .A2(n1280), .B1(A[49]), .B2(n1273), .ZN(n96) );
  AOI22_X1 U343 ( .A1(C[48]), .A2(n1277), .B1(A[48]), .B2(n1273), .ZN(n100) );
  AOI22_X1 U344 ( .A1(C[47]), .A2(n1279), .B1(A[47]), .B2(n1273), .ZN(n104) );
  AOI22_X1 U345 ( .A1(C[46]), .A2(n1280), .B1(A[46]), .B2(n1273), .ZN(n108) );
  AOI22_X1 U346 ( .A1(C[45]), .A2(n1277), .B1(A[45]), .B2(n1273), .ZN(n112) );
  AOI22_X1 U347 ( .A1(C[44]), .A2(n1281), .B1(A[44]), .B2(n1273), .ZN(n116) );
  AOI22_X1 U348 ( .A1(C[43]), .A2(n1276), .B1(A[43]), .B2(n1273), .ZN(n120) );
  AOI22_X1 U349 ( .A1(C[4]), .A2(n1278), .B1(A[4]), .B2(n1273), .ZN(n92) );
  NAND4_X1 U350 ( .A1(n260), .A2(n261), .A3(n262), .A4(n263), .ZN(Y[11]) );
  AOI22_X1 U351 ( .A1(G[11]), .A2(n1300), .B1(E[11]), .B2(n1294), .ZN(n262) );
  NAND4_X1 U352 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(Y[7]) );
  AOI22_X1 U353 ( .A1(F[7]), .A2(n1292), .B1(D[7]), .B2(n1286), .ZN(n29) );
  AOI22_X1 U354 ( .A1(G[7]), .A2(n1302), .B1(E[7]), .B2(n1298), .ZN(n30) );
  AOI22_X1 U355 ( .A1(G[10]), .A2(n1302), .B1(E[10]), .B2(n1299), .ZN(n6) );
  NOR3_X1 U356 ( .A1(n1319), .A2(SEL[1]), .A3(n1317), .ZN(n12) );
  NAND4_X1 U357 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(Y[3]) );
  NOR3_X1 U358 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1319), .ZN(n8) );
  INV_X1 U359 ( .A(SEL[1]), .ZN(n1318) );
  AOI22_X1 U360 ( .A1(C[42]), .A2(n1279), .B1(A[42]), .B2(n1272), .ZN(n124) );
  AOI22_X1 U361 ( .A1(C[41]), .A2(n1280), .B1(A[41]), .B2(n1272), .ZN(n128) );
  AOI22_X1 U362 ( .A1(C[40]), .A2(n1277), .B1(A[40]), .B2(n1272), .ZN(n132) );
  AOI22_X1 U363 ( .A1(C[39]), .A2(n1281), .B1(A[39]), .B2(n1272), .ZN(n140) );
  AOI22_X1 U364 ( .A1(C[36]), .A2(n1280), .B1(A[36]), .B2(n1272), .ZN(n152) );
  AOI22_X1 U365 ( .A1(C[37]), .A2(n1279), .B1(A[37]), .B2(n1272), .ZN(n148) );
  AOI22_X1 U366 ( .A1(C[38]), .A2(n1276), .B1(A[38]), .B2(n1272), .ZN(n144) );
  AOI22_X1 U367 ( .A1(C[35]), .A2(n1281), .B1(A[35]), .B2(n1272), .ZN(n156) );
  AOI22_X1 U368 ( .A1(C[32]), .A2(n1276), .B1(A[32]), .B2(n1272), .ZN(n168) );
  AOI22_X1 U369 ( .A1(C[34]), .A2(n1277), .B1(A[34]), .B2(n1272), .ZN(n160) );
  AOI22_X1 U370 ( .A1(C[33]), .A2(n1279), .B1(A[33]), .B2(n1272), .ZN(n164) );
  AOI22_X1 U371 ( .A1(C[3]), .A2(n1278), .B1(A[3]), .B2(n1272), .ZN(n136) );
  NOR3_X1 U372 ( .A1(n1319), .A2(SEL[2]), .A3(n1266), .ZN(n13) );
  NOR3_X1 U373 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n15) );
  INV_X1 U374 ( .A(SEL[2]), .ZN(n1317) );
  NAND4_X1 U375 ( .A1(n144), .A2(n145), .A3(n146), .A4(n147), .ZN(Y[38]) );
  AOI22_X1 U376 ( .A1(C[2]), .A2(n1279), .B1(A[2]), .B2(n1271), .ZN(n180) );
  CLKBUF_X3 U377 ( .A(n1269), .Z(n1277) );
  CLKBUF_X1 U378 ( .A(n15), .Z(n1275) );
  CLKBUF_X1 U379 ( .A(n1269), .Z(n1281) );
  CLKBUF_X1 U380 ( .A(n13), .Z(n1287) );
  CLKBUF_X1 U381 ( .A(n12), .Z(n1293) );
  CLKBUF_X1 U382 ( .A(n11), .Z(n1299) );
  CLKBUF_X1 U383 ( .A(n9), .Z(n1310) );
  CLKBUF_X1 U384 ( .A(n1265), .Z(n1316) );
endmodule


module MUX81_GENERIC_NBIT64_15 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382;

  NOR3_X2 U318 ( .A1(n1381), .A2(SEL[0]), .A3(n1380), .ZN(n9) );
  BUF_X1 U1 ( .A(n11), .Z(n1362) );
  BUF_X2 U2 ( .A(n1333), .Z(n1377) );
  INV_X1 U3 ( .A(n1381), .ZN(n1332) );
  BUF_X2 U4 ( .A(n1333), .Z(n1376) );
  CLKBUF_X2 U5 ( .A(n1333), .Z(n1378) );
  CLKBUF_X3 U6 ( .A(n1373), .Z(n1371) );
  BUF_X2 U7 ( .A(n9), .Z(n1373) );
  CLKBUF_X3 U8 ( .A(n9), .Z(n1370) );
  CLKBUF_X3 U9 ( .A(n1333), .Z(n1374) );
  BUF_X2 U10 ( .A(n12), .Z(n1355) );
  BUF_X1 U11 ( .A(n12), .Z(n1356) );
  BUF_X1 U12 ( .A(n12), .Z(n1354) );
  CLKBUF_X3 U13 ( .A(n11), .Z(n1361) );
  BUF_X1 U14 ( .A(n11), .Z(n1360) );
  NOR3_X2 U15 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1382), .ZN(n11) );
  AOI22_X1 U16 ( .A1(C[37]), .A2(n1377), .B1(G[37]), .B2(n1371), .ZN(n159) );
  AOI22_X1 U17 ( .A1(C[36]), .A2(n1378), .B1(G[36]), .B2(n1371), .ZN(n163) );
  AOI22_X1 U18 ( .A1(C[40]), .A2(n1379), .B1(G[40]), .B2(n1371), .ZN(n143) );
  AOI22_X1 U19 ( .A1(C[42]), .A2(n1374), .B1(G[42]), .B2(n1371), .ZN(n135) );
  AOI22_X1 U20 ( .A1(C[38]), .A2(n1374), .B1(G[38]), .B2(n1371), .ZN(n155) );
  BUF_X1 U21 ( .A(n15), .Z(n1335) );
  BUF_X1 U22 ( .A(n15), .Z(n1336) );
  BUF_X1 U23 ( .A(n15), .Z(n1337) );
  BUF_X1 U24 ( .A(n15), .Z(n1334) );
  BUF_X1 U25 ( .A(n15), .Z(n1338) );
  CLKBUF_X1 U26 ( .A(n11), .Z(n1359) );
  CLKBUF_X1 U27 ( .A(n11), .Z(n1358) );
  CLKBUF_X1 U28 ( .A(n1333), .Z(n1375) );
  CLKBUF_X1 U29 ( .A(n12), .Z(n1352) );
  CLKBUF_X1 U30 ( .A(n12), .Z(n1353) );
  BUF_X2 U31 ( .A(n9), .Z(n1372) );
  BUF_X1 U32 ( .A(n10), .Z(n1365) );
  BUF_X1 U33 ( .A(n14), .Z(n1341) );
  BUF_X1 U34 ( .A(n10), .Z(n1366) );
  BUF_X1 U35 ( .A(n14), .Z(n1342) );
  BUF_X1 U36 ( .A(n10), .Z(n1367) );
  BUF_X1 U37 ( .A(n14), .Z(n1343) );
  BUF_X1 U38 ( .A(n10), .Z(n1364) );
  BUF_X1 U39 ( .A(n14), .Z(n1340) );
  BUF_X1 U40 ( .A(n10), .Z(n1368) );
  BUF_X1 U41 ( .A(n14), .Z(n1344) );
  BUF_X1 U42 ( .A(n13), .Z(n1350) );
  BUF_X1 U43 ( .A(n13), .Z(n1349) );
  BUF_X1 U44 ( .A(n13), .Z(n1348) );
  BUF_X1 U45 ( .A(n13), .Z(n1346) );
  BUF_X1 U46 ( .A(n13), .Z(n1347) );
  AOI22_X1 U47 ( .A1(C[14]), .A2(n1374), .B1(G[14]), .B2(n1373), .ZN(n19) );
  AOI22_X1 U48 ( .A1(C[20]), .A2(n1377), .B1(G[20]), .B2(n1370), .ZN(n231) );
  AOI22_X1 U49 ( .A1(C[34]), .A2(n1375), .B1(G[34]), .B2(n1371), .ZN(n171) );
  AOI22_X1 U50 ( .A1(C[24]), .A2(n1374), .B1(G[24]), .B2(n1371), .ZN(n215) );
  INV_X1 U51 ( .A(SEL[0]), .ZN(n1382) );
  AOI22_X1 U52 ( .A1(C[25]), .A2(n1378), .B1(G[25]), .B2(n1371), .ZN(n211) );
  AOI22_X1 U53 ( .A1(C[9]), .A2(n1377), .B1(G[9]), .B2(n1373), .ZN(n27) );
  AOI22_X1 U54 ( .A1(C[21]), .A2(n1375), .B1(G[21]), .B2(n1370), .ZN(n227) );
  AOI22_X1 U55 ( .A1(C[28]), .A2(n1377), .B1(G[28]), .B2(n1371), .ZN(n199) );
  AOI22_X1 U56 ( .A1(C[10]), .A2(n1378), .B1(G[10]), .B2(n1370), .ZN(n263) );
  AOI22_X1 U57 ( .A1(C[11]), .A2(n1379), .B1(G[11]), .B2(n1370), .ZN(n259) );
  AOI22_X1 U58 ( .A1(C[29]), .A2(n1374), .B1(G[29]), .B2(n1371), .ZN(n195) );
  AOI22_X1 U59 ( .A1(C[26]), .A2(n1377), .B1(G[26]), .B2(n1371), .ZN(n207) );
  AOI22_X1 U60 ( .A1(C[30]), .A2(n1378), .B1(G[30]), .B2(n1371), .ZN(n187) );
  AOI22_X1 U61 ( .A1(A[4]), .A2(n1343), .B1(H[4]), .B2(n1337), .ZN(n100) );
  AOI22_X1 U62 ( .A1(E[4]), .A2(n1355), .B1(D[4]), .B2(n1349), .ZN(n101) );
  AOI22_X1 U63 ( .A1(F[4]), .A2(n1367), .B1(B[4]), .B2(n1362), .ZN(n102) );
  AOI22_X1 U64 ( .A1(E[12]), .A2(n1352), .B1(D[12]), .B2(n1346), .ZN(n253) );
  NAND4_X1 U65 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(Y[8]) );
  AOI22_X1 U66 ( .A1(A[8]), .A2(n1344), .B1(H[8]), .B2(n1338), .ZN(n28) );
  AOI22_X1 U67 ( .A1(E[8]), .A2(n1357), .B1(D[8]), .B2(n1350), .ZN(n29) );
  AOI22_X1 U68 ( .A1(F[8]), .A2(n1368), .B1(B[8]), .B2(n1361), .ZN(n30) );
  NAND4_X1 U69 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(Y[2]) );
  AOI22_X1 U70 ( .A1(A[2]), .A2(n1341), .B1(H[2]), .B2(n1335), .ZN(n188) );
  AOI22_X1 U71 ( .A1(C[2]), .A2(n1377), .B1(G[2]), .B2(n1371), .ZN(n191) );
  AOI22_X1 U72 ( .A1(E[2]), .A2(n1355), .B1(D[2]), .B2(n1347), .ZN(n189) );
  AOI22_X1 U73 ( .A1(A[15]), .A2(n1345), .B1(H[15]), .B2(n1339), .ZN(n4) );
  AOI22_X1 U74 ( .A1(F[15]), .A2(n1369), .B1(B[15]), .B2(n1361), .ZN(n6) );
  AOI22_X1 U75 ( .A1(C[15]), .A2(n1377), .B1(G[15]), .B2(n1373), .ZN(n7) );
  AOI22_X1 U76 ( .A1(A[22]), .A2(n1340), .B1(H[22]), .B2(n1334), .ZN(n220) );
  AOI22_X1 U77 ( .A1(F[22]), .A2(n1364), .B1(B[22]), .B2(n1360), .ZN(n222) );
  AOI22_X1 U78 ( .A1(A[33]), .A2(n1341), .B1(H[33]), .B2(n1335), .ZN(n172) );
  AOI22_X1 U79 ( .A1(F[33]), .A2(n1365), .B1(B[33]), .B2(n1361), .ZN(n174) );
  AOI22_X1 U80 ( .A1(C[33]), .A2(n1378), .B1(G[33]), .B2(n1371), .ZN(n175) );
  AOI22_X1 U81 ( .A1(A[30]), .A2(n1341), .B1(H[30]), .B2(n1335), .ZN(n184) );
  AOI22_X1 U82 ( .A1(F[30]), .A2(n1365), .B1(B[30]), .B2(n1361), .ZN(n186) );
  AOI22_X1 U83 ( .A1(A[3]), .A2(n1342), .B1(H[3]), .B2(n1336), .ZN(n144) );
  AOI22_X1 U84 ( .A1(E[3]), .A2(n1355), .B1(D[3]), .B2(n1348), .ZN(n145) );
  AOI22_X1 U85 ( .A1(F[3]), .A2(n1366), .B1(B[3]), .B2(n1362), .ZN(n146) );
  AOI22_X1 U86 ( .A1(A[23]), .A2(n1341), .B1(H[23]), .B2(n1335), .ZN(n216) );
  AOI22_X1 U87 ( .A1(F[23]), .A2(n1365), .B1(B[23]), .B2(n1361), .ZN(n218) );
  AOI22_X1 U88 ( .A1(E[23]), .A2(n1353), .B1(D[23]), .B2(n1347), .ZN(n217) );
  AOI22_X1 U89 ( .A1(A[5]), .A2(n1344), .B1(H[5]), .B2(n1338), .ZN(n56) );
  AOI22_X1 U90 ( .A1(E[5]), .A2(n1355), .B1(D[5]), .B2(n1350), .ZN(n57) );
  AOI22_X1 U91 ( .A1(A[38]), .A2(n1342), .B1(H[38]), .B2(n1336), .ZN(n152) );
  AOI22_X1 U92 ( .A1(F[38]), .A2(n1366), .B1(B[38]), .B2(n1360), .ZN(n154) );
  AOI22_X1 U93 ( .A1(E[38]), .A2(n1354), .B1(D[38]), .B2(n1348), .ZN(n153) );
  AOI22_X1 U94 ( .A1(A[19]), .A2(n1340), .B1(H[19]), .B2(n1334), .ZN(n236) );
  AOI22_X1 U95 ( .A1(F[19]), .A2(n1364), .B1(B[19]), .B2(n1358), .ZN(n238) );
  AOI22_X1 U96 ( .A1(C[19]), .A2(n1374), .B1(G[19]), .B2(n1370), .ZN(n239) );
  AOI22_X1 U97 ( .A1(E[48]), .A2(n1353), .B1(D[48]), .B2(n1349), .ZN(n109) );
  AOI22_X1 U98 ( .A1(E[52]), .A2(n1354), .B1(D[52]), .B2(n1349), .ZN(n89) );
  AOI22_X1 U99 ( .A1(E[53]), .A2(n1356), .B1(D[53]), .B2(n1349), .ZN(n85) );
  AOI22_X1 U100 ( .A1(E[50]), .A2(n1354), .B1(D[50]), .B2(n1349), .ZN(n97) );
  AOI22_X1 U101 ( .A1(E[45]), .A2(n1354), .B1(D[45]), .B2(n1349), .ZN(n121) );
  AOI22_X1 U102 ( .A1(E[46]), .A2(n1356), .B1(D[46]), .B2(n1349), .ZN(n117) );
  AOI22_X1 U103 ( .A1(E[54]), .A2(n1353), .B1(D[54]), .B2(n1349), .ZN(n81) );
  AOI22_X1 U104 ( .A1(E[51]), .A2(n1356), .B1(D[51]), .B2(n1349), .ZN(n93) );
  AOI22_X1 U105 ( .A1(E[47]), .A2(n1352), .B1(D[47]), .B2(n1349), .ZN(n113) );
  AOI22_X1 U106 ( .A1(E[55]), .A2(n1352), .B1(D[55]), .B2(n1349), .ZN(n77) );
  AOI22_X1 U107 ( .A1(E[56]), .A2(n1357), .B1(D[56]), .B2(n1350), .ZN(n73) );
  AOI22_X1 U108 ( .A1(E[57]), .A2(n1354), .B1(D[57]), .B2(n1350), .ZN(n69) );
  AOI22_X1 U109 ( .A1(E[63]), .A2(n1354), .B1(D[63]), .B2(n1350), .ZN(n41) );
  AOI22_X1 U110 ( .A1(E[61]), .A2(n1357), .B1(D[61]), .B2(n1350), .ZN(n49) );
  AOI22_X1 U111 ( .A1(E[62]), .A2(n1354), .B1(D[62]), .B2(n1350), .ZN(n45) );
  AOI22_X1 U112 ( .A1(E[59]), .A2(n1356), .B1(D[59]), .B2(n1350), .ZN(n61) );
  AOI22_X1 U113 ( .A1(E[58]), .A2(n1352), .B1(D[58]), .B2(n1350), .ZN(n65) );
  AOI22_X1 U114 ( .A1(E[60]), .A2(n1353), .B1(D[60]), .B2(n1350), .ZN(n53) );
  AOI22_X1 U115 ( .A1(E[41]), .A2(n1357), .B1(D[41]), .B2(n1348), .ZN(n137) );
  AOI22_X1 U116 ( .A1(E[44]), .A2(n1357), .B1(D[44]), .B2(n1348), .ZN(n125) );
  AOI22_X1 U117 ( .A1(A[35]), .A2(n1342), .B1(H[35]), .B2(n1336), .ZN(n164) );
  AOI22_X1 U118 ( .A1(F[35]), .A2(n1366), .B1(B[35]), .B2(n1363), .ZN(n166) );
  AOI22_X1 U119 ( .A1(A[16]), .A2(n1340), .B1(H[16]), .B2(n1334), .ZN(n248) );
  AOI22_X1 U120 ( .A1(F[16]), .A2(n1364), .B1(B[16]), .B2(n1359), .ZN(n250) );
  AOI22_X1 U121 ( .A1(A[17]), .A2(n1340), .B1(H[17]), .B2(n1334), .ZN(n244) );
  AOI22_X1 U122 ( .A1(F[17]), .A2(n1364), .B1(B[17]), .B2(n1360), .ZN(n246) );
  AOI22_X1 U123 ( .A1(A[31]), .A2(n1341), .B1(H[31]), .B2(n1335), .ZN(n180) );
  AOI22_X1 U124 ( .A1(F[31]), .A2(n1365), .B1(B[31]), .B2(n1361), .ZN(n182) );
  AOI22_X1 U125 ( .A1(A[27]), .A2(n1341), .B1(H[27]), .B2(n1335), .ZN(n200) );
  AOI22_X1 U126 ( .A1(F[27]), .A2(n1365), .B1(B[27]), .B2(n1359), .ZN(n202) );
  AOI22_X1 U127 ( .A1(A[43]), .A2(n1342), .B1(H[43]), .B2(n1336), .ZN(n128) );
  AOI22_X1 U128 ( .A1(F[43]), .A2(n1366), .B1(B[43]), .B2(n1361), .ZN(n130) );
  AOI22_X1 U129 ( .A1(E[43]), .A2(n1353), .B1(D[43]), .B2(n1348), .ZN(n129) );
  AOI22_X1 U130 ( .A1(E[13]), .A2(n1357), .B1(D[13]), .B2(n1351), .ZN(n21) );
  AOI22_X1 U131 ( .A1(E[32]), .A2(n1354), .B1(D[32]), .B2(n1347), .ZN(n177) );
  AOI22_X1 U132 ( .A1(F[2]), .A2(n1365), .B1(B[2]), .B2(n1362), .ZN(n190) );
  NAND4_X1 U133 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(Y[7]) );
  AOI22_X1 U134 ( .A1(A[7]), .A2(n1344), .B1(H[7]), .B2(n1338), .ZN(n32) );
  AOI22_X1 U135 ( .A1(E[7]), .A2(n1355), .B1(D[7]), .B2(n1350), .ZN(n33) );
  AOI22_X1 U136 ( .A1(F[7]), .A2(n1368), .B1(B[7]), .B2(n1362), .ZN(n34) );
  NAND4_X1 U137 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(Y[13]) );
  AOI22_X1 U138 ( .A1(A[13]), .A2(n1345), .B1(H[13]), .B2(n1339), .ZN(n20) );
  AOI22_X1 U139 ( .A1(F[13]), .A2(n1369), .B1(B[13]), .B2(n1361), .ZN(n22) );
  AOI22_X1 U140 ( .A1(C[13]), .A2(n1378), .B1(G[13]), .B2(n1373), .ZN(n23) );
  AOI22_X1 U141 ( .A1(A[29]), .A2(n1341), .B1(H[29]), .B2(n1335), .ZN(n192) );
  AOI22_X1 U142 ( .A1(F[29]), .A2(n1365), .B1(B[29]), .B2(n1363), .ZN(n194) );
  AOI22_X1 U143 ( .A1(A[26]), .A2(n1341), .B1(H[26]), .B2(n1335), .ZN(n204) );
  AOI22_X1 U144 ( .A1(F[26]), .A2(n1365), .B1(B[26]), .B2(n1360), .ZN(n206) );
  AOI22_X1 U145 ( .A1(E[39]), .A2(n1352), .B1(D[39]), .B2(n1348), .ZN(n149) );
  AOI22_X1 U146 ( .A1(A[39]), .A2(n1342), .B1(H[39]), .B2(n1336), .ZN(n148) );
  AOI22_X1 U147 ( .A1(F[39]), .A2(n1366), .B1(B[39]), .B2(n1359), .ZN(n150) );
  AOI22_X1 U148 ( .A1(C[39]), .A2(n1375), .B1(G[39]), .B2(n1371), .ZN(n151) );
  NAND4_X1 U149 ( .A1(n240), .A2(n241), .A3(n242), .A4(n243), .ZN(Y[18]) );
  AOI22_X1 U150 ( .A1(A[18]), .A2(n1340), .B1(H[18]), .B2(n1334), .ZN(n240) );
  AOI22_X1 U151 ( .A1(F[18]), .A2(n1364), .B1(B[18]), .B2(n1363), .ZN(n242) );
  AOI22_X1 U152 ( .A1(C[18]), .A2(n1378), .B1(G[18]), .B2(n1370), .ZN(n243) );
  AOI22_X1 U153 ( .A1(E[49]), .A2(n1357), .B1(D[49]), .B2(n1349), .ZN(n105) );
  AOI22_X1 U154 ( .A1(E[19]), .A2(n1357), .B1(D[19]), .B2(n1346), .ZN(n237) );
  NAND4_X1 U155 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(Y[6]) );
  AOI22_X1 U156 ( .A1(A[6]), .A2(n1344), .B1(H[6]), .B2(n1338), .ZN(n36) );
  AOI22_X1 U157 ( .A1(E[6]), .A2(n1355), .B1(D[6]), .B2(n1350), .ZN(n37) );
  AOI22_X1 U158 ( .A1(F[6]), .A2(n1368), .B1(B[6]), .B2(n1362), .ZN(n38) );
  NAND4_X1 U159 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(Y[56]) );
  AOI22_X1 U160 ( .A1(A[56]), .A2(n1344), .B1(H[56]), .B2(n1338), .ZN(n72) );
  AOI22_X1 U161 ( .A1(F[56]), .A2(n1368), .B1(B[56]), .B2(n1363), .ZN(n74) );
  NAND4_X1 U162 ( .A1(n68), .A2(n69), .A3(n70), .A4(n71), .ZN(Y[57]) );
  AOI22_X1 U163 ( .A1(A[57]), .A2(n1344), .B1(H[57]), .B2(n1338), .ZN(n68) );
  AOI22_X1 U164 ( .A1(F[57]), .A2(n1368), .B1(B[57]), .B2(n1358), .ZN(n70) );
  NAND4_X1 U165 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(Y[58]) );
  AOI22_X1 U166 ( .A1(A[58]), .A2(n1344), .B1(H[58]), .B2(n1338), .ZN(n64) );
  AOI22_X1 U167 ( .A1(F[58]), .A2(n1368), .B1(B[58]), .B2(n1359), .ZN(n66) );
  NAND4_X1 U168 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .ZN(Y[61]) );
  AOI22_X1 U169 ( .A1(A[61]), .A2(n1344), .B1(H[61]), .B2(n1338), .ZN(n48) );
  AOI22_X1 U170 ( .A1(F[61]), .A2(n1368), .B1(B[61]), .B2(n1358), .ZN(n50) );
  NAND4_X1 U171 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(Y[62]) );
  AOI22_X1 U172 ( .A1(A[62]), .A2(n1344), .B1(H[62]), .B2(n1338), .ZN(n44) );
  AOI22_X1 U173 ( .A1(F[62]), .A2(n1368), .B1(B[62]), .B2(n1360), .ZN(n46) );
  NAND4_X1 U174 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(Y[63]) );
  AOI22_X1 U175 ( .A1(A[63]), .A2(n1344), .B1(H[63]), .B2(n1338), .ZN(n40) );
  AOI22_X1 U176 ( .A1(F[63]), .A2(n1368), .B1(B[63]), .B2(n1360), .ZN(n42) );
  NAND4_X1 U177 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(Y[60]) );
  AOI22_X1 U178 ( .A1(A[60]), .A2(n1344), .B1(H[60]), .B2(n1338), .ZN(n52) );
  AOI22_X1 U179 ( .A1(F[60]), .A2(n1368), .B1(B[60]), .B2(n1363), .ZN(n54) );
  NAND4_X1 U180 ( .A1(n88), .A2(n89), .A3(n90), .A4(n91), .ZN(Y[52]) );
  AOI22_X1 U181 ( .A1(A[52]), .A2(n1343), .B1(H[52]), .B2(n1337), .ZN(n88) );
  AOI22_X1 U182 ( .A1(F[52]), .A2(n1367), .B1(B[52]), .B2(n1358), .ZN(n90) );
  NAND4_X1 U183 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(Y[48]) );
  AOI22_X1 U184 ( .A1(A[48]), .A2(n1343), .B1(H[48]), .B2(n1337), .ZN(n108) );
  AOI22_X1 U185 ( .A1(F[48]), .A2(n1367), .B1(B[48]), .B2(n1360), .ZN(n110) );
  NAND4_X1 U186 ( .A1(n84), .A2(n85), .A3(n86), .A4(n87), .ZN(Y[53]) );
  AOI22_X1 U187 ( .A1(A[53]), .A2(n1343), .B1(H[53]), .B2(n1337), .ZN(n84) );
  AOI22_X1 U188 ( .A1(F[53]), .A2(n1367), .B1(B[53]), .B2(n1361), .ZN(n86) );
  NAND4_X1 U189 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(Y[49]) );
  AOI22_X1 U190 ( .A1(A[49]), .A2(n1343), .B1(H[49]), .B2(n1337), .ZN(n104) );
  AOI22_X1 U191 ( .A1(F[49]), .A2(n1367), .B1(B[49]), .B2(n1361), .ZN(n106) );
  NAND4_X1 U192 ( .A1(n96), .A2(n97), .A3(n98), .A4(n99), .ZN(Y[50]) );
  AOI22_X1 U193 ( .A1(A[50]), .A2(n1343), .B1(H[50]), .B2(n1337), .ZN(n96) );
  AOI22_X1 U194 ( .A1(F[50]), .A2(n1367), .B1(B[50]), .B2(n1359), .ZN(n98) );
  NAND4_X1 U195 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(Y[54]) );
  AOI22_X1 U196 ( .A1(A[54]), .A2(n1343), .B1(H[54]), .B2(n1337), .ZN(n80) );
  AOI22_X1 U197 ( .A1(F[54]), .A2(n1367), .B1(B[54]), .B2(n1359), .ZN(n82) );
  NAND4_X1 U198 ( .A1(n120), .A2(n121), .A3(n122), .A4(n123), .ZN(Y[45]) );
  AOI22_X1 U199 ( .A1(A[45]), .A2(n1343), .B1(H[45]), .B2(n1337), .ZN(n120) );
  AOI22_X1 U200 ( .A1(F[45]), .A2(n1367), .B1(B[45]), .B2(n1363), .ZN(n122) );
  NAND4_X1 U201 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(Y[46]) );
  AOI22_X1 U202 ( .A1(A[46]), .A2(n1343), .B1(H[46]), .B2(n1337), .ZN(n116) );
  AOI22_X1 U203 ( .A1(F[46]), .A2(n1367), .B1(B[46]), .B2(n1358), .ZN(n118) );
  NAND4_X1 U204 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(Y[47]) );
  AOI22_X1 U205 ( .A1(A[47]), .A2(n1343), .B1(H[47]), .B2(n1337), .ZN(n112) );
  AOI22_X1 U206 ( .A1(F[47]), .A2(n1367), .B1(B[47]), .B2(n1361), .ZN(n114) );
  NAND4_X1 U207 ( .A1(n156), .A2(n157), .A3(n158), .A4(n159), .ZN(Y[37]) );
  AOI22_X1 U208 ( .A1(A[37]), .A2(n1342), .B1(H[37]), .B2(n1336), .ZN(n156) );
  AOI22_X1 U209 ( .A1(F[37]), .A2(n1366), .B1(B[37]), .B2(n1361), .ZN(n158) );
  AOI22_X1 U210 ( .A1(E[37]), .A2(n1356), .B1(D[37]), .B2(n1348), .ZN(n157) );
  NAND4_X1 U211 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(Y[36]) );
  AOI22_X1 U212 ( .A1(A[36]), .A2(n1342), .B1(H[36]), .B2(n1336), .ZN(n160) );
  AOI22_X1 U213 ( .A1(F[36]), .A2(n1366), .B1(B[36]), .B2(n1358), .ZN(n162) );
  AOI22_X1 U214 ( .A1(E[36]), .A2(n1357), .B1(D[36]), .B2(n1348), .ZN(n161) );
  NAND4_X1 U215 ( .A1(n168), .A2(n169), .A3(n170), .A4(n171), .ZN(Y[34]) );
  AOI22_X1 U216 ( .A1(A[34]), .A2(n1342), .B1(H[34]), .B2(n1336), .ZN(n168) );
  AOI22_X1 U217 ( .A1(F[34]), .A2(n1366), .B1(B[34]), .B2(n1359), .ZN(n170) );
  AOI22_X1 U218 ( .A1(E[34]), .A2(n1352), .B1(D[34]), .B2(n1348), .ZN(n169) );
  NAND4_X1 U219 ( .A1(n140), .A2(n141), .A3(n142), .A4(n143), .ZN(Y[40]) );
  AOI22_X1 U220 ( .A1(A[40]), .A2(n1342), .B1(H[40]), .B2(n1336), .ZN(n140) );
  AOI22_X1 U221 ( .A1(F[40]), .A2(n1366), .B1(B[40]), .B2(n1363), .ZN(n142) );
  AOI22_X1 U222 ( .A1(E[40]), .A2(n1353), .B1(D[40]), .B2(n1348), .ZN(n141) );
  NAND4_X1 U223 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(Y[41]) );
  AOI22_X1 U224 ( .A1(A[41]), .A2(n1342), .B1(H[41]), .B2(n1336), .ZN(n136) );
  AOI22_X1 U225 ( .A1(F[41]), .A2(n1366), .B1(B[41]), .B2(n1358), .ZN(n138) );
  AOI22_X1 U226 ( .A1(C[41]), .A2(n1378), .B1(G[41]), .B2(n1371), .ZN(n139) );
  NAND4_X1 U227 ( .A1(n124), .A2(n125), .A3(n126), .A4(n127), .ZN(Y[44]) );
  AOI22_X1 U228 ( .A1(A[44]), .A2(n1342), .B1(H[44]), .B2(n1336), .ZN(n124) );
  AOI22_X1 U229 ( .A1(F[44]), .A2(n1366), .B1(B[44]), .B2(n1359), .ZN(n126) );
  AOI22_X1 U230 ( .A1(C[44]), .A2(n1375), .B1(G[44]), .B2(n1371), .ZN(n127) );
  NAND4_X1 U231 ( .A1(n132), .A2(n133), .A3(n134), .A4(n135), .ZN(Y[42]) );
  AOI22_X1 U232 ( .A1(A[42]), .A2(n1342), .B1(H[42]), .B2(n1336), .ZN(n132) );
  AOI22_X1 U233 ( .A1(F[42]), .A2(n1366), .B1(B[42]), .B2(n1360), .ZN(n134) );
  AOI22_X1 U234 ( .A1(E[42]), .A2(n1352), .B1(D[42]), .B2(n1348), .ZN(n133) );
  NAND4_X1 U235 ( .A1(n260), .A2(n261), .A3(n262), .A4(n263), .ZN(Y[10]) );
  AOI22_X1 U236 ( .A1(A[10]), .A2(n1340), .B1(H[10]), .B2(n1334), .ZN(n260) );
  AOI22_X1 U237 ( .A1(F[10]), .A2(n1364), .B1(B[10]), .B2(n1358), .ZN(n262) );
  AOI22_X1 U238 ( .A1(E[10]), .A2(n1353), .B1(D[10]), .B2(n1346), .ZN(n261) );
  NAND4_X1 U239 ( .A1(n228), .A2(n229), .A3(n230), .A4(n231), .ZN(Y[20]) );
  AOI22_X1 U240 ( .A1(A[20]), .A2(n1340), .B1(H[20]), .B2(n1334), .ZN(n228) );
  AOI22_X1 U241 ( .A1(F[20]), .A2(n1364), .B1(B[20]), .B2(n1361), .ZN(n230) );
  AOI22_X1 U242 ( .A1(E[20]), .A2(n1354), .B1(D[20]), .B2(n1346), .ZN(n229) );
  NAND4_X1 U243 ( .A1(n224), .A2(n225), .A3(n226), .A4(n227), .ZN(Y[21]) );
  AOI22_X1 U244 ( .A1(A[21]), .A2(n1340), .B1(H[21]), .B2(n1334), .ZN(n224) );
  AOI22_X1 U245 ( .A1(F[21]), .A2(n1364), .B1(B[21]), .B2(n1361), .ZN(n226) );
  AOI22_X1 U246 ( .A1(E[21]), .A2(n1356), .B1(D[21]), .B2(n1346), .ZN(n225) );
  NAND4_X1 U247 ( .A1(n252), .A2(n253), .A3(n254), .A4(n255), .ZN(Y[12]) );
  AOI22_X1 U248 ( .A1(A[12]), .A2(n1340), .B1(H[12]), .B2(n1334), .ZN(n252) );
  AOI22_X1 U249 ( .A1(F[12]), .A2(n1364), .B1(B[12]), .B2(n1358), .ZN(n254) );
  AOI22_X1 U250 ( .A1(C[12]), .A2(n1378), .B1(G[12]), .B2(n1370), .ZN(n255) );
  NAND4_X1 U251 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(Y[11]) );
  AOI22_X1 U252 ( .A1(A[11]), .A2(n1340), .B1(H[11]), .B2(n1334), .ZN(n256) );
  AOI22_X1 U253 ( .A1(F[11]), .A2(n1364), .B1(B[11]), .B2(n1359), .ZN(n258) );
  AOI22_X1 U254 ( .A1(E[11]), .A2(n1356), .B1(D[11]), .B2(n1346), .ZN(n257) );
  NAND4_X1 U255 ( .A1(n27), .A2(n25), .A3(n26), .A4(n24), .ZN(Y[9]) );
  AOI22_X1 U256 ( .A1(A[9]), .A2(n1345), .B1(H[9]), .B2(n1339), .ZN(n24) );
  AOI22_X1 U257 ( .A1(E[9]), .A2(n1354), .B1(D[9]), .B2(n1351), .ZN(n25) );
  AOI22_X1 U258 ( .A1(F[9]), .A2(n1369), .B1(B[9]), .B2(n1360), .ZN(n26) );
  NAND4_X1 U259 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(Y[14]) );
  AOI22_X1 U260 ( .A1(A[14]), .A2(n1345), .B1(H[14]), .B2(n1339), .ZN(n16) );
  AOI22_X1 U261 ( .A1(F[14]), .A2(n1369), .B1(B[14]), .B2(n1363), .ZN(n18) );
  AOI22_X1 U262 ( .A1(E[14]), .A2(n1353), .B1(D[14]), .B2(n1351), .ZN(n17) );
  NAND4_X1 U263 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(Y[32]) );
  AOI22_X1 U264 ( .A1(A[32]), .A2(n1341), .B1(H[32]), .B2(n1335), .ZN(n176) );
  AOI22_X1 U265 ( .A1(F[32]), .A2(n1365), .B1(B[32]), .B2(n1361), .ZN(n178) );
  AOI22_X1 U266 ( .A1(C[32]), .A2(n1377), .B1(G[32]), .B2(n1371), .ZN(n179) );
  NAND4_X1 U267 ( .A1(n212), .A2(n213), .A3(n214), .A4(n215), .ZN(Y[24]) );
  AOI22_X1 U268 ( .A1(A[24]), .A2(n1341), .B1(H[24]), .B2(n1335), .ZN(n212) );
  AOI22_X1 U269 ( .A1(F[24]), .A2(n1365), .B1(B[24]), .B2(n1361), .ZN(n214) );
  AOI22_X1 U270 ( .A1(E[24]), .A2(n1354), .B1(D[24]), .B2(n1347), .ZN(n213) );
  NAND4_X1 U271 ( .A1(n196), .A2(n197), .A3(n198), .A4(n199), .ZN(Y[28]) );
  AOI22_X1 U272 ( .A1(A[28]), .A2(n1341), .B1(H[28]), .B2(n1335), .ZN(n196) );
  AOI22_X1 U273 ( .A1(F[28]), .A2(n1365), .B1(B[28]), .B2(n1358), .ZN(n198) );
  AOI22_X1 U274 ( .A1(E[28]), .A2(n1352), .B1(D[28]), .B2(n1347), .ZN(n197) );
  NAND4_X1 U275 ( .A1(n208), .A2(n209), .A3(n210), .A4(n211), .ZN(Y[25]) );
  AOI22_X1 U276 ( .A1(A[25]), .A2(n1341), .B1(H[25]), .B2(n1335), .ZN(n208) );
  AOI22_X1 U277 ( .A1(F[25]), .A2(n1365), .B1(B[25]), .B2(n1361), .ZN(n210) );
  AOI22_X1 U278 ( .A1(E[25]), .A2(n1356), .B1(D[25]), .B2(n1347), .ZN(n209) );
  AOI22_X1 U279 ( .A1(F[5]), .A2(n1368), .B1(B[5]), .B2(n1362), .ZN(n58) );
  NAND4_X1 U280 ( .A1(n60), .A2(n61), .A3(n62), .A4(n63), .ZN(Y[59]) );
  AOI22_X1 U281 ( .A1(A[59]), .A2(n1344), .B1(H[59]), .B2(n1338), .ZN(n60) );
  AOI22_X1 U282 ( .A1(F[59]), .A2(n1368), .B1(B[59]), .B2(n1360), .ZN(n62) );
  NAND4_X1 U283 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(Y[51]) );
  AOI22_X1 U284 ( .A1(A[51]), .A2(n1343), .B1(H[51]), .B2(n1337), .ZN(n92) );
  AOI22_X1 U285 ( .A1(F[51]), .A2(n1367), .B1(B[51]), .B2(n1363), .ZN(n94) );
  NAND4_X1 U286 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(Y[55]) );
  AOI22_X1 U287 ( .A1(A[55]), .A2(n1343), .B1(H[55]), .B2(n1337), .ZN(n76) );
  AOI22_X1 U288 ( .A1(F[55]), .A2(n1367), .B1(B[55]), .B2(n1360), .ZN(n78) );
  NAND4_X1 U289 ( .A1(n232), .A2(n233), .A3(n234), .A4(n235), .ZN(Y[1]) );
  AOI22_X1 U290 ( .A1(A[1]), .A2(n1340), .B1(H[1]), .B2(n1334), .ZN(n232) );
  AOI22_X1 U291 ( .A1(F[1]), .A2(n1364), .B1(B[1]), .B2(n1361), .ZN(n234) );
  AOI22_X1 U292 ( .A1(E[1]), .A2(n1356), .B1(D[1]), .B2(n1346), .ZN(n233) );
  NAND4_X1 U293 ( .A1(n264), .A2(n265), .A3(n266), .A4(n267), .ZN(Y[0]) );
  AOI22_X1 U294 ( .A1(A[0]), .A2(n1340), .B1(H[0]), .B2(n1334), .ZN(n264) );
  AOI22_X1 U295 ( .A1(E[0]), .A2(n1356), .B1(D[0]), .B2(n1346), .ZN(n265) );
  AOI22_X1 U296 ( .A1(F[0]), .A2(n1364), .B1(B[0]), .B2(n1361), .ZN(n266) );
  AOI22_X1 U297 ( .A1(C[1]), .A2(n1377), .B1(G[1]), .B2(n1370), .ZN(n235) );
  AOI22_X1 U298 ( .A1(C[0]), .A2(n1377), .B1(G[0]), .B2(n1370), .ZN(n267) );
  NAND4_X1 U299 ( .A1(n100), .A2(n101), .A3(n102), .A4(n103), .ZN(Y[4]) );
  BUF_X2 U300 ( .A(n8), .Z(n1333) );
  NOR3_X1 U301 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1381), .ZN(n8) );
  AOI22_X1 U302 ( .A1(E[27]), .A2(n1354), .B1(D[27]), .B2(n1347), .ZN(n201) );
  NAND4_X1 U303 ( .A1(n236), .A2(n237), .A3(n238), .A4(n239), .ZN(Y[19]) );
  NAND4_X1 U304 ( .A1(n221), .A2(n220), .A3(n222), .A4(n223), .ZN(Y[22]) );
  AOI22_X1 U305 ( .A1(E[17]), .A2(n1356), .B1(D[17]), .B2(n1346), .ZN(n245) );
  AOI22_X1 U306 ( .A1(E[16]), .A2(n1352), .B1(D[16]), .B2(n1346), .ZN(n249) );
  AOI22_X1 U307 ( .A1(C[17]), .A2(n1377), .B1(G[17]), .B2(n1370), .ZN(n247) );
  NAND4_X1 U308 ( .A1(n144), .A2(n145), .A3(n146), .A4(n147), .ZN(Y[3]) );
  AOI22_X1 U309 ( .A1(C[22]), .A2(n1379), .B1(G[22]), .B2(n1370), .ZN(n223) );
  AOI22_X1 U310 ( .A1(E[18]), .A2(n1353), .B1(D[18]), .B2(n1346), .ZN(n241) );
  AOI22_X1 U311 ( .A1(C[27]), .A2(n1378), .B1(G[27]), .B2(n1371), .ZN(n203) );
  AOI22_X1 U312 ( .A1(E[35]), .A2(n1353), .B1(D[35]), .B2(n1348), .ZN(n165) );
  NAND4_X1 U313 ( .A1(n248), .A2(n249), .A3(n250), .A4(n251), .ZN(Y[16]) );
  NAND4_X1 U314 ( .A1(n184), .A2(n185), .A3(n186), .A4(n187), .ZN(Y[30]) );
  AOI22_X1 U315 ( .A1(E[30]), .A2(n1353), .B1(D[30]), .B2(n1347), .ZN(n185) );
  AOI22_X1 U316 ( .A1(E[22]), .A2(n1352), .B1(D[22]), .B2(n1346), .ZN(n221) );
  AOI22_X1 U317 ( .A1(E[31]), .A2(n1357), .B1(D[31]), .B2(n1347), .ZN(n181) );
  AOI22_X1 U319 ( .A1(C[31]), .A2(n1374), .B1(G[31]), .B2(n1371), .ZN(n183) );
  AOI22_X1 U320 ( .A1(C[3]), .A2(n1376), .B1(G[3]), .B2(n1373), .ZN(n147) );
  NOR3_X1 U321 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n15) );
  NAND4_X1 U322 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(Y[43]) );
  NAND4_X1 U323 ( .A1(n192), .A2(n193), .A3(n194), .A4(n195), .ZN(Y[29]) );
  NAND4_X1 U324 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(Y[33]) );
  AOI22_X1 U325 ( .A1(C[63]), .A2(n1374), .B1(G[63]), .B2(n1371), .ZN(n43) );
  AOI22_X1 U326 ( .A1(C[62]), .A2(n1379), .B1(G[62]), .B2(n1371), .ZN(n47) );
  AOI22_X1 U327 ( .A1(C[61]), .A2(n1375), .B1(G[61]), .B2(n1371), .ZN(n51) );
  AOI22_X1 U328 ( .A1(C[60]), .A2(n1378), .B1(G[60]), .B2(n1371), .ZN(n55) );
  AOI22_X1 U329 ( .A1(C[58]), .A2(n1374), .B1(G[58]), .B2(n1371), .ZN(n67) );
  AOI22_X1 U330 ( .A1(C[59]), .A2(n1379), .B1(G[59]), .B2(n1371), .ZN(n63) );
  AOI22_X1 U331 ( .A1(C[57]), .A2(n1375), .B1(G[57]), .B2(n1371), .ZN(n71) );
  AOI22_X1 U332 ( .A1(C[56]), .A2(n1378), .B1(G[56]), .B2(n1371), .ZN(n75) );
  AOI22_X1 U333 ( .A1(C[8]), .A2(n1375), .B1(G[8]), .B2(n1370), .ZN(n31) );
  NAND4_X1 U334 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(Y[5]) );
  AOI22_X1 U335 ( .A1(C[7]), .A2(n1376), .B1(G[7]), .B2(n1370), .ZN(n35) );
  AOI22_X1 U336 ( .A1(C[6]), .A2(n1376), .B1(G[6]), .B2(n1373), .ZN(n39) );
  AOI22_X1 U337 ( .A1(C[5]), .A2(n1376), .B1(G[5]), .B2(n1373), .ZN(n59) );
  NAND4_X1 U338 ( .A1(n204), .A2(n205), .A3(n206), .A4(n207), .ZN(Y[26]) );
  AOI22_X1 U339 ( .A1(E[26]), .A2(n1357), .B1(D[26]), .B2(n1347), .ZN(n205) );
  AOI22_X1 U340 ( .A1(E[15]), .A2(n1354), .B1(D[15]), .B2(n1351), .ZN(n5) );
  AOI22_X1 U341 ( .A1(C[16]), .A2(n1374), .B1(G[16]), .B2(n1370), .ZN(n251) );
  AOI22_X1 U342 ( .A1(C[43]), .A2(n1377), .B1(G[43]), .B2(n1371), .ZN(n131) );
  AOI22_X1 U343 ( .A1(E[33]), .A2(n1356), .B1(D[33]), .B2(n1347), .ZN(n173) );
  AOI22_X1 U344 ( .A1(C[23]), .A2(n1378), .B1(G[23]), .B2(n1371), .ZN(n219) );
  NAND4_X1 U345 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(Y[27]) );
  AOI22_X1 U346 ( .A1(E[29]), .A2(n1356), .B1(D[29]), .B2(n1347), .ZN(n193) );
  NOR3_X1 U347 ( .A1(n1380), .A2(n1332), .A3(n1382), .ZN(n10) );
  AOI22_X1 U348 ( .A1(C[54]), .A2(n1374), .B1(G[54]), .B2(n1372), .ZN(n83) );
  AOI22_X1 U349 ( .A1(C[55]), .A2(n1378), .B1(G[55]), .B2(n1372), .ZN(n79) );
  AOI22_X1 U350 ( .A1(C[53]), .A2(n1377), .B1(G[53]), .B2(n1372), .ZN(n87) );
  AOI22_X1 U351 ( .A1(C[52]), .A2(n1374), .B1(G[52]), .B2(n1372), .ZN(n91) );
  AOI22_X1 U352 ( .A1(C[51]), .A2(n1379), .B1(G[51]), .B2(n1372), .ZN(n95) );
  AOI22_X1 U353 ( .A1(C[50]), .A2(n1375), .B1(G[50]), .B2(n1372), .ZN(n99) );
  AOI22_X1 U354 ( .A1(C[49]), .A2(n1378), .B1(G[49]), .B2(n1372), .ZN(n107) );
  AOI22_X1 U355 ( .A1(C[48]), .A2(n1377), .B1(G[48]), .B2(n1372), .ZN(n111) );
  AOI22_X1 U356 ( .A1(C[47]), .A2(n1374), .B1(G[47]), .B2(n1372), .ZN(n115) );
  AOI22_X1 U357 ( .A1(C[46]), .A2(n1378), .B1(G[46]), .B2(n1372), .ZN(n119) );
  AOI22_X1 U358 ( .A1(C[45]), .A2(n1379), .B1(G[45]), .B2(n1372), .ZN(n123) );
  AOI22_X1 U359 ( .A1(C[4]), .A2(n1376), .B1(G[4]), .B2(n1372), .ZN(n103) );
  NOR3_X1 U360 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1380), .ZN(n12) );
  INV_X1 U361 ( .A(SEL[1]), .ZN(n1381) );
  NAND4_X1 U362 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(Y[15]) );
  NAND4_X1 U363 ( .A1(n244), .A2(n245), .A3(n246), .A4(n247), .ZN(Y[17]) );
  AOI22_X1 U364 ( .A1(C[35]), .A2(n1379), .B1(G[35]), .B2(n1371), .ZN(n167) );
  NOR3_X1 U365 ( .A1(n1381), .A2(SEL[2]), .A3(n1382), .ZN(n13) );
  NOR3_X1 U366 ( .A1(n1332), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  INV_X1 U367 ( .A(SEL[2]), .ZN(n1380) );
  NAND4_X1 U368 ( .A1(n148), .A2(n149), .A3(n150), .A4(n151), .ZN(Y[39]) );
  NAND4_X1 U369 ( .A1(n216), .A2(n217), .A3(n218), .A4(n219), .ZN(Y[23]) );
  NAND4_X1 U370 ( .A1(n152), .A2(n153), .A3(n154), .A4(n155), .ZN(Y[38]) );
  NAND4_X1 U371 ( .A1(n180), .A2(n181), .A3(n182), .A4(n183), .ZN(Y[31]) );
  NAND4_X1 U372 ( .A1(n164), .A2(n165), .A3(n166), .A4(n167), .ZN(Y[35]) );
  CLKBUF_X1 U373 ( .A(n15), .Z(n1339) );
  CLKBUF_X1 U374 ( .A(n14), .Z(n1345) );
  CLKBUF_X1 U375 ( .A(n13), .Z(n1351) );
  CLKBUF_X1 U376 ( .A(n12), .Z(n1357) );
  CLKBUF_X1 U377 ( .A(n11), .Z(n1363) );
  CLKBUF_X1 U378 ( .A(n10), .Z(n1369) );
  CLKBUF_X1 U379 ( .A(n1333), .Z(n1379) );
endmodule


module MUX81_GENERIC_NBIT64_14 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455;

  NAND4_X1 U1 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AND3_X1 U2 ( .A1(SEL[1]), .A2(n1455), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U3 ( .A1(n190), .A2(n188), .A3(n187), .ZN(n1405) );
  NAND2_X1 U4 ( .A1(n189), .A2(n1405), .ZN(Y[27]) );
  CLKBUF_X1 U5 ( .A(n12), .Z(n1421) );
  BUF_X2 U6 ( .A(n12), .Z(n1422) );
  CLKBUF_X1 U7 ( .A(n12), .Z(n1419) );
  CLKBUF_X1 U8 ( .A(n12), .Z(n1420) );
  BUF_X2 U9 ( .A(n10), .Z(n1433) );
  BUF_X2 U10 ( .A(n10), .Z(n1434) );
  CLKBUF_X1 U11 ( .A(n10), .Z(n1431) );
  CLKBUF_X1 U12 ( .A(n10), .Z(n1432) );
  BUF_X1 U13 ( .A(n13), .Z(n1415) );
  BUF_X1 U14 ( .A(n13), .Z(n1413) );
  BUF_X1 U15 ( .A(n13), .Z(n1412) );
  BUF_X1 U16 ( .A(n13), .Z(n1416) );
  BUF_X1 U17 ( .A(n13), .Z(n1414) );
  BUF_X1 U18 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U19 ( .A(n8), .Z(n1443) );
  CLKBUF_X1 U20 ( .A(n8), .Z(n1442) );
  BUF_X1 U21 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U22 ( .A(n8), .Z(n1446) );
  CLKBUF_X1 U23 ( .A(n8), .Z(n1444) );
  CLKBUF_X1 U24 ( .A(n8), .Z(n1445) );
  BUF_X1 U25 ( .A(n11), .Z(n1427) );
  BUF_X1 U26 ( .A(n11), .Z(n1425) );
  BUF_X1 U27 ( .A(n11), .Z(n1426) );
  BUF_X1 U28 ( .A(n11), .Z(n1424) );
  BUF_X1 U29 ( .A(n11), .Z(n1428) );
  BUF_X1 U30 ( .A(n7), .Z(n1448) );
  BUF_X1 U31 ( .A(n7), .Z(n1449) );
  BUF_X1 U32 ( .A(n7), .Z(n1450) );
  BUF_X1 U33 ( .A(n9), .Z(n1439) );
  BUF_X1 U34 ( .A(n7), .Z(n1451) );
  BUF_X1 U35 ( .A(n9), .Z(n1440) );
  BUF_X1 U36 ( .A(n9), .Z(n1437) );
  BUF_X1 U37 ( .A(n9), .Z(n1438) );
  BUF_X1 U38 ( .A(n9), .Z(n1436) );
  BUF_X1 U39 ( .A(n7), .Z(n1452) );
  BUF_X1 U40 ( .A(n14), .Z(n1409) );
  BUF_X1 U41 ( .A(n14), .Z(n1407) );
  BUF_X1 U42 ( .A(n14), .Z(n1408) );
  BUF_X1 U43 ( .A(n14), .Z(n1406) );
  BUF_X1 U44 ( .A(n14), .Z(n1410) );
  NOR3_X1 U45 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1455), .ZN(n13) );
  NOR3_X1 U46 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1454), .ZN(n12) );
  AND3_X1 U47 ( .A1(n1455), .A2(n1454), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U48 ( .A(SEL[1]), .ZN(n1454) );
  INV_X1 U49 ( .A(SEL[0]), .ZN(n1455) );
  NOR3_X1 U50 ( .A1(n1455), .A2(SEL[2]), .A3(n1454), .ZN(n11) );
  NOR3_X1 U51 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U52 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U53 ( .A1(SEL[0]), .A2(n1454), .A3(SEL[2]), .ZN(n9) );
  AOI22_X1 U54 ( .A1(H[6]), .A2(n1453), .B1(G[6]), .B2(n1447), .ZN(n26) );
  AOI22_X1 U55 ( .A1(B[6]), .A2(n1417), .B1(A[6]), .B2(n1411), .ZN(n23) );
  AOI22_X1 U56 ( .A1(D[6]), .A2(n1429), .B1(C[6]), .B2(n1423), .ZN(n24) );
  AOI22_X1 U57 ( .A1(F[44]), .A2(n1439), .B1(E[44]), .B2(n1433), .ZN(n113) );
  AOI22_X1 U58 ( .A1(F[42]), .A2(n1439), .B1(E[42]), .B2(n1433), .ZN(n121) );
  AOI22_X1 U59 ( .A1(F[46]), .A2(n1439), .B1(E[46]), .B2(n1433), .ZN(n105) );
  AOI22_X1 U60 ( .A1(F[38]), .A2(n1438), .B1(E[38]), .B2(n1432), .ZN(n141) );
  AOI22_X1 U61 ( .A1(F[43]), .A2(n1439), .B1(E[43]), .B2(n1433), .ZN(n117) );
  AOI22_X1 U62 ( .A1(F[47]), .A2(n1439), .B1(E[47]), .B2(n1433), .ZN(n101) );
  AOI22_X1 U63 ( .A1(F[24]), .A2(n1437), .B1(E[24]), .B2(n1431), .ZN(n201) );
  NAND4_X1 U64 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U65 ( .A1(B[15]), .A2(n1412), .B1(A[15]), .B2(n1406), .ZN(n239) );
  AOI22_X1 U66 ( .A1(D[15]), .A2(n1424), .B1(C[15]), .B2(n1418), .ZN(n240) );
  AOI22_X1 U67 ( .A1(H[15]), .A2(n1448), .B1(G[15]), .B2(n1442), .ZN(n242) );
  NAND4_X1 U68 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U69 ( .A1(H[8]), .A2(n1453), .B1(G[8]), .B2(n1447), .ZN(n18) );
  AOI22_X1 U70 ( .A1(B[8]), .A2(n1417), .B1(A[8]), .B2(n1411), .ZN(n15) );
  AOI22_X1 U71 ( .A1(D[8]), .A2(n1429), .B1(C[8]), .B2(n1423), .ZN(n16) );
  AOI22_X1 U72 ( .A1(H[10]), .A2(n1448), .B1(G[10]), .B2(n1442), .ZN(n262) );
  AOI22_X1 U73 ( .A1(H[11]), .A2(n1448), .B1(G[11]), .B2(n1442), .ZN(n258) );
  AOI22_X1 U74 ( .A1(H[9]), .A2(n1453), .B1(G[9]), .B2(n1447), .ZN(n6) );
  NAND4_X1 U75 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U76 ( .A1(D[4]), .A2(n1427), .B1(C[4]), .B2(n1421), .ZN(n88) );
  AOI22_X1 U77 ( .A1(H[4]), .A2(n1451), .B1(G[4]), .B2(n1445), .ZN(n90) );
  AOI22_X1 U78 ( .A1(B[4]), .A2(n1415), .B1(A[4]), .B2(n1409), .ZN(n87) );
  NAND4_X1 U79 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U80 ( .A1(B[9]), .A2(n1417), .B1(A[9]), .B2(n1411), .ZN(n3) );
  AOI22_X1 U81 ( .A1(F[9]), .A2(n1441), .B1(E[9]), .B2(n1435), .ZN(n5) );
  AOI22_X1 U82 ( .A1(D[9]), .A2(n1429), .B1(C[9]), .B2(n1423), .ZN(n4) );
  AOI22_X1 U83 ( .A1(F[33]), .A2(n1438), .B1(E[33]), .B2(n1432), .ZN(n161) );
  AOI22_X1 U84 ( .A1(F[36]), .A2(n1438), .B1(E[36]), .B2(n1432), .ZN(n149) );
  AOI22_X1 U85 ( .A1(F[40]), .A2(n1438), .B1(E[40]), .B2(n1432), .ZN(n129) );
  AOI22_X1 U86 ( .A1(F[32]), .A2(n1438), .B1(E[32]), .B2(n1432), .ZN(n165) );
  AOI22_X1 U87 ( .A1(F[34]), .A2(n1438), .B1(E[34]), .B2(n1432), .ZN(n157) );
  AOI22_X1 U88 ( .A1(F[52]), .A2(n1439), .B1(E[52]), .B2(n1433), .ZN(n77) );
  AOI22_X1 U89 ( .A1(F[18]), .A2(n1436), .B1(E[18]), .B2(n1430), .ZN(n229) );
  AOI22_X1 U90 ( .A1(F[35]), .A2(n1438), .B1(E[35]), .B2(n1432), .ZN(n153) );
  AOI22_X1 U91 ( .A1(F[48]), .A2(n1439), .B1(E[48]), .B2(n1433), .ZN(n97) );
  AOI22_X1 U92 ( .A1(F[19]), .A2(n1436), .B1(E[19]), .B2(n1430), .ZN(n225) );
  AOI22_X1 U93 ( .A1(F[49]), .A2(n1439), .B1(E[49]), .B2(n1433), .ZN(n93) );
  AOI22_X1 U94 ( .A1(F[20]), .A2(n1437), .B1(E[20]), .B2(n1431), .ZN(n217) );
  AOI22_X1 U95 ( .A1(F[50]), .A2(n1439), .B1(E[50]), .B2(n1433), .ZN(n85) );
  AOI22_X1 U96 ( .A1(F[28]), .A2(n1437), .B1(E[28]), .B2(n1431), .ZN(n185) );
  AOI22_X1 U97 ( .A1(F[21]), .A2(n1437), .B1(E[21]), .B2(n1431), .ZN(n213) );
  AOI22_X1 U98 ( .A1(F[53]), .A2(n1440), .B1(E[53]), .B2(n1434), .ZN(n73) );
  AOI22_X1 U99 ( .A1(F[39]), .A2(n1438), .B1(E[39]), .B2(n1432), .ZN(n137) );
  AOI22_X1 U100 ( .A1(F[54]), .A2(n1440), .B1(E[54]), .B2(n1434), .ZN(n69) );
  AOI22_X1 U101 ( .A1(F[25]), .A2(n1437), .B1(E[25]), .B2(n1431), .ZN(n197) );
  AOI22_X1 U102 ( .A1(F[26]), .A2(n1437), .B1(E[26]), .B2(n1431), .ZN(n193) );
  AOI22_X1 U103 ( .A1(F[30]), .A2(n1437), .B1(E[30]), .B2(n1431), .ZN(n173) );
  AOI22_X1 U104 ( .A1(F[27]), .A2(n1437), .B1(E[27]), .B2(n1431), .ZN(n189) );
  AOI22_X1 U105 ( .A1(F[51]), .A2(n1439), .B1(E[51]), .B2(n1433), .ZN(n81) );
  AOI22_X1 U106 ( .A1(F[4]), .A2(n1439), .B1(E[4]), .B2(n1433), .ZN(n89) );
  AOI22_X1 U107 ( .A1(F[22]), .A2(n1437), .B1(E[22]), .B2(n1431), .ZN(n209) );
  AOI22_X1 U108 ( .A1(F[13]), .A2(n1436), .B1(E[13]), .B2(n1430), .ZN(n249) );
  AOI22_X1 U109 ( .A1(F[14]), .A2(n1436), .B1(E[14]), .B2(n1430), .ZN(n245) );
  AOI22_X1 U110 ( .A1(F[23]), .A2(n1437), .B1(E[23]), .B2(n1431), .ZN(n205) );
  AOI22_X1 U111 ( .A1(F[15]), .A2(n1436), .B1(E[15]), .B2(n1430), .ZN(n241) );
  AOI22_X1 U112 ( .A1(F[12]), .A2(n1436), .B1(E[12]), .B2(n1430), .ZN(n253) );
  AOI22_X1 U113 ( .A1(F[55]), .A2(n1440), .B1(E[55]), .B2(n1434), .ZN(n65) );
  AOI22_X1 U114 ( .A1(F[56]), .A2(n1440), .B1(E[56]), .B2(n1434), .ZN(n61) );
  AOI22_X1 U115 ( .A1(F[57]), .A2(n1440), .B1(E[57]), .B2(n1434), .ZN(n57) );
  AOI22_X1 U116 ( .A1(F[58]), .A2(n1440), .B1(E[58]), .B2(n1434), .ZN(n53) );
  AOI22_X1 U117 ( .A1(F[60]), .A2(n1440), .B1(E[60]), .B2(n1434), .ZN(n41) );
  AOI22_X1 U118 ( .A1(F[5]), .A2(n1440), .B1(E[5]), .B2(n1434), .ZN(n45) );
  AOI22_X1 U119 ( .A1(F[59]), .A2(n1440), .B1(E[59]), .B2(n1434), .ZN(n49) );
  AOI22_X1 U120 ( .A1(F[61]), .A2(n1440), .B1(E[61]), .B2(n1434), .ZN(n37) );
  AOI22_X1 U121 ( .A1(F[62]), .A2(n1440), .B1(E[62]), .B2(n1434), .ZN(n33) );
  AOI22_X1 U122 ( .A1(F[63]), .A2(n1440), .B1(E[63]), .B2(n1434), .ZN(n29) );
  AOI22_X1 U123 ( .A1(F[6]), .A2(n1441), .B1(E[6]), .B2(n1435), .ZN(n25) );
  AOI22_X1 U124 ( .A1(F[8]), .A2(n1441), .B1(E[8]), .B2(n1435), .ZN(n17) );
  NAND4_X1 U125 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U126 ( .A1(B[13]), .A2(n1412), .B1(A[13]), .B2(n1406), .ZN(n247) );
  AOI22_X1 U127 ( .A1(H[13]), .A2(n1448), .B1(G[13]), .B2(n1442), .ZN(n250) );
  AOI22_X1 U128 ( .A1(D[13]), .A2(n1424), .B1(C[13]), .B2(n1418), .ZN(n248) );
  AOI22_X1 U129 ( .A1(D[7]), .A2(n1429), .B1(C[7]), .B2(n1423), .ZN(n20) );
  NAND4_X1 U130 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U131 ( .A1(B[10]), .A2(n1412), .B1(A[10]), .B2(n1406), .ZN(n259) );
  AOI22_X1 U132 ( .A1(D[10]), .A2(n1424), .B1(C[10]), .B2(n1418), .ZN(n260) );
  AOI22_X1 U133 ( .A1(F[10]), .A2(n1436), .B1(E[10]), .B2(n1430), .ZN(n261) );
  NAND4_X1 U134 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U135 ( .A1(B[12]), .A2(n1412), .B1(A[12]), .B2(n1406), .ZN(n251) );
  AOI22_X1 U136 ( .A1(H[12]), .A2(n1448), .B1(G[12]), .B2(n1442), .ZN(n254) );
  AOI22_X1 U137 ( .A1(D[12]), .A2(n1424), .B1(C[12]), .B2(n1418), .ZN(n252) );
  NAND4_X1 U138 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U139 ( .A1(B[22]), .A2(n1413), .B1(A[22]), .B2(n1407), .ZN(n207) );
  AOI22_X1 U140 ( .A1(D[22]), .A2(n1425), .B1(C[22]), .B2(n1419), .ZN(n208) );
  AOI22_X1 U141 ( .A1(H[22]), .A2(n1449), .B1(G[22]), .B2(n1443), .ZN(n210) );
  NAND4_X1 U142 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U143 ( .A1(B[11]), .A2(n1412), .B1(A[11]), .B2(n1406), .ZN(n255) );
  AOI22_X1 U144 ( .A1(D[11]), .A2(n1424), .B1(C[11]), .B2(n1418), .ZN(n256) );
  AOI22_X1 U145 ( .A1(F[11]), .A2(n1436), .B1(E[11]), .B2(n1430), .ZN(n257) );
  NAND4_X1 U146 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U147 ( .A1(H[5]), .A2(n1452), .B1(G[5]), .B2(n1446), .ZN(n46) );
  AOI22_X1 U148 ( .A1(B[5]), .A2(n1416), .B1(A[5]), .B2(n1410), .ZN(n43) );
  AOI22_X1 U149 ( .A1(D[5]), .A2(n1428), .B1(C[5]), .B2(n1422), .ZN(n44) );
  NAND4_X1 U150 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U151 ( .A1(B[33]), .A2(n1414), .B1(A[33]), .B2(n1408), .ZN(n159) );
  AOI22_X1 U152 ( .A1(D[33]), .A2(n1426), .B1(C[33]), .B2(n1420), .ZN(n160) );
  AOI22_X1 U153 ( .A1(H[33]), .A2(n1450), .B1(G[33]), .B2(n1444), .ZN(n162) );
  NAND4_X1 U154 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U155 ( .A1(B[37]), .A2(n1414), .B1(A[37]), .B2(n1408), .ZN(n143) );
  AOI22_X1 U156 ( .A1(D[37]), .A2(n1426), .B1(C[37]), .B2(n1420), .ZN(n144) );
  AOI22_X1 U157 ( .A1(H[37]), .A2(n1450), .B1(G[37]), .B2(n1444), .ZN(n146) );
  NAND4_X1 U158 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U159 ( .A1(B[20]), .A2(n1413), .B1(A[20]), .B2(n1407), .ZN(n215) );
  AOI22_X1 U160 ( .A1(D[20]), .A2(n1425), .B1(C[20]), .B2(n1419), .ZN(n216) );
  AOI22_X1 U161 ( .A1(H[20]), .A2(n1449), .B1(G[20]), .B2(n1443), .ZN(n218) );
  NAND4_X1 U162 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U163 ( .A1(B[32]), .A2(n1414), .B1(A[32]), .B2(n1408), .ZN(n163) );
  AOI22_X1 U164 ( .A1(D[32]), .A2(n1426), .B1(C[32]), .B2(n1420), .ZN(n164) );
  AOI22_X1 U165 ( .A1(H[32]), .A2(n1450), .B1(G[32]), .B2(n1444), .ZN(n166) );
  NAND4_X1 U166 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U167 ( .A1(B[36]), .A2(n1414), .B1(A[36]), .B2(n1408), .ZN(n147) );
  AOI22_X1 U168 ( .A1(D[36]), .A2(n1426), .B1(C[36]), .B2(n1420), .ZN(n148) );
  AOI22_X1 U169 ( .A1(H[36]), .A2(n1450), .B1(G[36]), .B2(n1444), .ZN(n150) );
  NAND4_X1 U170 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U171 ( .A1(B[29]), .A2(n1413), .B1(A[29]), .B2(n1407), .ZN(n179) );
  AOI22_X1 U172 ( .A1(D[29]), .A2(n1425), .B1(C[29]), .B2(n1419), .ZN(n180) );
  AOI22_X1 U173 ( .A1(H[29]), .A2(n1449), .B1(G[29]), .B2(n1443), .ZN(n182) );
  NAND4_X1 U174 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U175 ( .A1(B[16]), .A2(n1412), .B1(A[16]), .B2(n1406), .ZN(n235) );
  AOI22_X1 U176 ( .A1(H[16]), .A2(n1448), .B1(G[16]), .B2(n1442), .ZN(n238) );
  AOI22_X1 U177 ( .A1(D[16]), .A2(n1424), .B1(C[16]), .B2(n1418), .ZN(n236) );
  NAND4_X1 U178 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U179 ( .A1(B[40]), .A2(n1414), .B1(A[40]), .B2(n1408), .ZN(n127) );
  AOI22_X1 U180 ( .A1(D[40]), .A2(n1426), .B1(C[40]), .B2(n1420), .ZN(n128) );
  AOI22_X1 U181 ( .A1(H[40]), .A2(n1450), .B1(G[40]), .B2(n1444), .ZN(n130) );
  NAND4_X1 U182 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U183 ( .A1(B[52]), .A2(n1415), .B1(A[52]), .B2(n1409), .ZN(n75) );
  AOI22_X1 U184 ( .A1(D[52]), .A2(n1427), .B1(C[52]), .B2(n1421), .ZN(n76) );
  AOI22_X1 U185 ( .A1(H[52]), .A2(n1451), .B1(G[52]), .B2(n1445), .ZN(n78) );
  NAND4_X1 U186 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U187 ( .A1(B[21]), .A2(n1413), .B1(A[21]), .B2(n1407), .ZN(n211) );
  AOI22_X1 U188 ( .A1(D[21]), .A2(n1425), .B1(C[21]), .B2(n1419), .ZN(n212) );
  AOI22_X1 U189 ( .A1(H[21]), .A2(n1449), .B1(G[21]), .B2(n1443), .ZN(n214) );
  NAND4_X1 U190 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U191 ( .A1(B[53]), .A2(n1416), .B1(A[53]), .B2(n1410), .ZN(n71) );
  AOI22_X1 U192 ( .A1(D[53]), .A2(n1428), .B1(C[53]), .B2(n1422), .ZN(n72) );
  AOI22_X1 U193 ( .A1(H[53]), .A2(n1452), .B1(G[53]), .B2(n1446), .ZN(n74) );
  NAND4_X1 U194 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U195 ( .A1(B[17]), .A2(n1412), .B1(A[17]), .B2(n1406), .ZN(n231) );
  AOI22_X1 U196 ( .A1(D[17]), .A2(n1424), .B1(C[17]), .B2(n1418), .ZN(n232) );
  AOI22_X1 U197 ( .A1(H[17]), .A2(n1448), .B1(G[17]), .B2(n1442), .ZN(n234) );
  NAND4_X1 U198 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U199 ( .A1(B[24]), .A2(n1413), .B1(A[24]), .B2(n1407), .ZN(n199) );
  AOI22_X1 U200 ( .A1(D[24]), .A2(n1425), .B1(C[24]), .B2(n1419), .ZN(n200) );
  AOI22_X1 U201 ( .A1(H[24]), .A2(n1449), .B1(G[24]), .B2(n1443), .ZN(n202) );
  NAND4_X1 U202 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U203 ( .A1(B[48]), .A2(n1415), .B1(A[48]), .B2(n1409), .ZN(n95) );
  AOI22_X1 U204 ( .A1(D[48]), .A2(n1427), .B1(C[48]), .B2(n1421), .ZN(n96) );
  AOI22_X1 U205 ( .A1(H[48]), .A2(n1451), .B1(G[48]), .B2(n1445), .ZN(n98) );
  NAND4_X1 U206 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U207 ( .A1(B[54]), .A2(n1416), .B1(A[54]), .B2(n1410), .ZN(n67) );
  AOI22_X1 U208 ( .A1(D[54]), .A2(n1428), .B1(C[54]), .B2(n1422), .ZN(n68) );
  AOI22_X1 U209 ( .A1(H[54]), .A2(n1452), .B1(G[54]), .B2(n1446), .ZN(n70) );
  NAND4_X1 U210 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U211 ( .A1(B[38]), .A2(n1414), .B1(A[38]), .B2(n1408), .ZN(n139) );
  AOI22_X1 U212 ( .A1(D[38]), .A2(n1426), .B1(C[38]), .B2(n1420), .ZN(n140) );
  AOI22_X1 U213 ( .A1(H[38]), .A2(n1450), .B1(G[38]), .B2(n1444), .ZN(n142) );
  NAND4_X1 U214 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U215 ( .A1(B[34]), .A2(n1414), .B1(A[34]), .B2(n1408), .ZN(n155) );
  AOI22_X1 U216 ( .A1(D[34]), .A2(n1426), .B1(C[34]), .B2(n1420), .ZN(n156) );
  AOI22_X1 U217 ( .A1(H[34]), .A2(n1450), .B1(G[34]), .B2(n1444), .ZN(n158) );
  NAND4_X1 U218 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U219 ( .A1(B[28]), .A2(n1413), .B1(A[28]), .B2(n1407), .ZN(n183) );
  AOI22_X1 U220 ( .A1(D[28]), .A2(n1425), .B1(C[28]), .B2(n1419), .ZN(n184) );
  AOI22_X1 U221 ( .A1(H[28]), .A2(n1449), .B1(G[28]), .B2(n1443), .ZN(n186) );
  NAND4_X1 U222 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U223 ( .A1(B[49]), .A2(n1415), .B1(A[49]), .B2(n1409), .ZN(n91) );
  AOI22_X1 U224 ( .A1(D[49]), .A2(n1427), .B1(C[49]), .B2(n1421), .ZN(n92) );
  AOI22_X1 U225 ( .A1(H[49]), .A2(n1451), .B1(G[49]), .B2(n1445), .ZN(n94) );
  NAND4_X1 U226 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U227 ( .A1(B[41]), .A2(n1414), .B1(A[41]), .B2(n1408), .ZN(n123) );
  AOI22_X1 U228 ( .A1(D[41]), .A2(n1426), .B1(C[41]), .B2(n1420), .ZN(n124) );
  AOI22_X1 U229 ( .A1(H[41]), .A2(n1450), .B1(G[41]), .B2(n1444), .ZN(n126) );
  NAND4_X1 U230 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U231 ( .A1(B[26]), .A2(n1413), .B1(A[26]), .B2(n1407), .ZN(n191) );
  AOI22_X1 U232 ( .A1(D[26]), .A2(n1425), .B1(C[26]), .B2(n1419), .ZN(n192) );
  AOI22_X1 U233 ( .A1(H[26]), .A2(n1449), .B1(G[26]), .B2(n1443), .ZN(n194) );
  NAND4_X1 U234 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U235 ( .A1(B[44]), .A2(n1415), .B1(A[44]), .B2(n1409), .ZN(n111) );
  AOI22_X1 U236 ( .A1(D[44]), .A2(n1427), .B1(C[44]), .B2(n1421), .ZN(n112) );
  AOI22_X1 U237 ( .A1(H[44]), .A2(n1451), .B1(G[44]), .B2(n1445), .ZN(n114) );
  NAND4_X1 U238 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U239 ( .A1(B[50]), .A2(n1415), .B1(A[50]), .B2(n1409), .ZN(n83) );
  AOI22_X1 U240 ( .A1(D[50]), .A2(n1427), .B1(C[50]), .B2(n1421), .ZN(n84) );
  AOI22_X1 U241 ( .A1(H[50]), .A2(n1451), .B1(G[50]), .B2(n1445), .ZN(n86) );
  NAND4_X1 U242 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U243 ( .A1(B[30]), .A2(n1413), .B1(A[30]), .B2(n1407), .ZN(n171) );
  AOI22_X1 U244 ( .A1(D[30]), .A2(n1425), .B1(C[30]), .B2(n1419), .ZN(n172) );
  AOI22_X1 U245 ( .A1(H[30]), .A2(n1449), .B1(G[30]), .B2(n1443), .ZN(n174) );
  NAND4_X1 U246 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U247 ( .A1(B[45]), .A2(n1415), .B1(A[45]), .B2(n1409), .ZN(n107) );
  AOI22_X1 U248 ( .A1(D[45]), .A2(n1427), .B1(C[45]), .B2(n1421), .ZN(n108) );
  AOI22_X1 U249 ( .A1(H[45]), .A2(n1451), .B1(G[45]), .B2(n1445), .ZN(n110) );
  NAND4_X1 U250 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U251 ( .A1(B[42]), .A2(n1415), .B1(A[42]), .B2(n1409), .ZN(n119) );
  AOI22_X1 U252 ( .A1(D[42]), .A2(n1427), .B1(C[42]), .B2(n1421), .ZN(n120) );
  AOI22_X1 U253 ( .A1(H[42]), .A2(n1451), .B1(G[42]), .B2(n1445), .ZN(n122) );
  NAND4_X1 U254 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U255 ( .A1(B[14]), .A2(n1412), .B1(A[14]), .B2(n1406), .ZN(n243) );
  AOI22_X1 U256 ( .A1(D[14]), .A2(n1424), .B1(C[14]), .B2(n1418), .ZN(n244) );
  AOI22_X1 U257 ( .A1(H[14]), .A2(n1448), .B1(G[14]), .B2(n1442), .ZN(n246) );
  NAND4_X1 U258 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U259 ( .A1(B[46]), .A2(n1415), .B1(A[46]), .B2(n1409), .ZN(n103) );
  AOI22_X1 U260 ( .A1(D[46]), .A2(n1427), .B1(C[46]), .B2(n1421), .ZN(n104) );
  AOI22_X1 U261 ( .A1(H[46]), .A2(n1451), .B1(G[46]), .B2(n1445), .ZN(n106) );
  NAND4_X1 U262 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U263 ( .A1(B[51]), .A2(n1415), .B1(A[51]), .B2(n1409), .ZN(n79) );
  AOI22_X1 U264 ( .A1(D[51]), .A2(n1427), .B1(C[51]), .B2(n1421), .ZN(n80) );
  AOI22_X1 U265 ( .A1(H[51]), .A2(n1451), .B1(G[51]), .B2(n1445), .ZN(n82) );
  NAND4_X1 U266 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U267 ( .A1(B[56]), .A2(n1416), .B1(A[56]), .B2(n1410), .ZN(n59) );
  AOI22_X1 U268 ( .A1(D[56]), .A2(n1428), .B1(C[56]), .B2(n1422), .ZN(n60) );
  AOI22_X1 U269 ( .A1(H[56]), .A2(n1452), .B1(G[56]), .B2(n1446), .ZN(n62) );
  NAND4_X1 U270 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U271 ( .A1(B[57]), .A2(n1416), .B1(A[57]), .B2(n1410), .ZN(n55) );
  AOI22_X1 U272 ( .A1(D[57]), .A2(n1428), .B1(C[57]), .B2(n1422), .ZN(n56) );
  AOI22_X1 U273 ( .A1(H[57]), .A2(n1452), .B1(G[57]), .B2(n1446), .ZN(n58) );
  NAND4_X1 U274 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U275 ( .A1(B[58]), .A2(n1416), .B1(A[58]), .B2(n1410), .ZN(n51) );
  AOI22_X1 U276 ( .A1(D[58]), .A2(n1428), .B1(C[58]), .B2(n1422), .ZN(n52) );
  AOI22_X1 U277 ( .A1(H[58]), .A2(n1452), .B1(G[58]), .B2(n1446), .ZN(n54) );
  NAND4_X1 U278 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U279 ( .A1(B[60]), .A2(n1416), .B1(A[60]), .B2(n1410), .ZN(n39) );
  AOI22_X1 U280 ( .A1(D[60]), .A2(n1428), .B1(C[60]), .B2(n1422), .ZN(n40) );
  AOI22_X1 U281 ( .A1(H[60]), .A2(n1452), .B1(G[60]), .B2(n1446), .ZN(n42) );
  NAND4_X1 U282 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U283 ( .A1(B[61]), .A2(n1416), .B1(A[61]), .B2(n1410), .ZN(n35) );
  AOI22_X1 U284 ( .A1(D[61]), .A2(n1428), .B1(C[61]), .B2(n1422), .ZN(n36) );
  AOI22_X1 U285 ( .A1(H[61]), .A2(n1452), .B1(G[61]), .B2(n1446), .ZN(n38) );
  NAND4_X1 U286 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U287 ( .A1(B[62]), .A2(n1416), .B1(A[62]), .B2(n1410), .ZN(n31) );
  AOI22_X1 U288 ( .A1(D[62]), .A2(n1428), .B1(C[62]), .B2(n1422), .ZN(n32) );
  AOI22_X1 U289 ( .A1(H[62]), .A2(n1452), .B1(G[62]), .B2(n1446), .ZN(n34) );
  NAND4_X1 U290 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U291 ( .A1(B[63]), .A2(n1416), .B1(A[63]), .B2(n1410), .ZN(n27) );
  AOI22_X1 U292 ( .A1(D[63]), .A2(n1428), .B1(C[63]), .B2(n1422), .ZN(n28) );
  AOI22_X1 U293 ( .A1(H[63]), .A2(n1452), .B1(G[63]), .B2(n1446), .ZN(n30) );
  AOI22_X1 U294 ( .A1(F[41]), .A2(n1438), .B1(E[41]), .B2(n1432), .ZN(n125) );
  NAND4_X1 U295 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U296 ( .A1(B[19]), .A2(n1412), .B1(A[19]), .B2(n1406), .ZN(n223) );
  AOI22_X1 U297 ( .A1(D[19]), .A2(n1424), .B1(C[19]), .B2(n1418), .ZN(n224) );
  AOI22_X1 U298 ( .A1(H[19]), .A2(n1448), .B1(G[19]), .B2(n1442), .ZN(n226) );
  AOI22_X1 U299 ( .A1(F[17]), .A2(n1436), .B1(E[17]), .B2(n1430), .ZN(n233) );
  AOI22_X1 U300 ( .A1(F[45]), .A2(n1439), .B1(E[45]), .B2(n1433), .ZN(n109) );
  NAND4_X1 U301 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U302 ( .A1(B[55]), .A2(n1416), .B1(A[55]), .B2(n1410), .ZN(n63) );
  AOI22_X1 U303 ( .A1(D[55]), .A2(n1428), .B1(C[55]), .B2(n1422), .ZN(n64) );
  AOI22_X1 U304 ( .A1(H[55]), .A2(n1452), .B1(G[55]), .B2(n1446), .ZN(n66) );
  NAND4_X1 U305 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U306 ( .A1(B[59]), .A2(n1416), .B1(A[59]), .B2(n1410), .ZN(n47) );
  AOI22_X1 U307 ( .A1(D[59]), .A2(n1428), .B1(C[59]), .B2(n1422), .ZN(n48) );
  AOI22_X1 U308 ( .A1(H[59]), .A2(n1452), .B1(G[59]), .B2(n1446), .ZN(n50) );
  NAND4_X1 U309 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U310 ( .A1(B[23]), .A2(n1413), .B1(A[23]), .B2(n1407), .ZN(n203) );
  AOI22_X1 U311 ( .A1(D[23]), .A2(n1425), .B1(C[23]), .B2(n1419), .ZN(n204) );
  AOI22_X1 U312 ( .A1(H[23]), .A2(n1449), .B1(G[23]), .B2(n1443), .ZN(n206) );
  NAND4_X1 U313 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U314 ( .A1(B[18]), .A2(n1412), .B1(A[18]), .B2(n1406), .ZN(n227) );
  AOI22_X1 U315 ( .A1(D[18]), .A2(n1424), .B1(C[18]), .B2(n1418), .ZN(n228) );
  AOI22_X1 U316 ( .A1(H[18]), .A2(n1448), .B1(G[18]), .B2(n1442), .ZN(n230) );
  NAND4_X1 U317 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U318 ( .A1(B[25]), .A2(n1413), .B1(A[25]), .B2(n1407), .ZN(n195) );
  AOI22_X1 U319 ( .A1(D[25]), .A2(n1425), .B1(C[25]), .B2(n1419), .ZN(n196) );
  AOI22_X1 U320 ( .A1(H[25]), .A2(n1449), .B1(G[25]), .B2(n1443), .ZN(n198) );
  NAND4_X1 U321 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U322 ( .A1(B[39]), .A2(n1414), .B1(A[39]), .B2(n1408), .ZN(n135) );
  AOI22_X1 U323 ( .A1(D[39]), .A2(n1426), .B1(C[39]), .B2(n1420), .ZN(n136) );
  AOI22_X1 U324 ( .A1(H[39]), .A2(n1450), .B1(G[39]), .B2(n1444), .ZN(n138) );
  NAND4_X1 U325 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U326 ( .A1(B[43]), .A2(n1415), .B1(A[43]), .B2(n1409), .ZN(n115) );
  AOI22_X1 U327 ( .A1(D[43]), .A2(n1427), .B1(C[43]), .B2(n1421), .ZN(n116) );
  AOI22_X1 U328 ( .A1(H[43]), .A2(n1451), .B1(G[43]), .B2(n1445), .ZN(n118) );
  NAND4_X1 U329 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U330 ( .A1(B[47]), .A2(n1415), .B1(A[47]), .B2(n1409), .ZN(n99) );
  AOI22_X1 U331 ( .A1(D[47]), .A2(n1427), .B1(C[47]), .B2(n1421), .ZN(n100) );
  AOI22_X1 U332 ( .A1(H[47]), .A2(n1451), .B1(G[47]), .B2(n1445), .ZN(n102) );
  AOI22_X1 U333 ( .A1(F[29]), .A2(n1437), .B1(E[29]), .B2(n1431), .ZN(n181) );
  NAND4_X1 U334 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U335 ( .A1(H[7]), .A2(n1453), .B1(G[7]), .B2(n1447), .ZN(n22) );
  AOI22_X1 U336 ( .A1(B[7]), .A2(n1417), .B1(A[7]), .B2(n1411), .ZN(n19) );
  AOI22_X1 U337 ( .A1(F[7]), .A2(n1441), .B1(E[7]), .B2(n1435), .ZN(n21) );
  NAND4_X1 U338 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U339 ( .A1(B[31]), .A2(n1414), .B1(A[31]), .B2(n1408), .ZN(n167) );
  AOI22_X1 U340 ( .A1(D[31]), .A2(n1426), .B1(C[31]), .B2(n1420), .ZN(n168) );
  AOI22_X1 U341 ( .A1(H[31]), .A2(n1450), .B1(G[31]), .B2(n1444), .ZN(n170) );
  AOI22_X1 U342 ( .A1(F[16]), .A2(n1436), .B1(E[16]), .B2(n1430), .ZN(n237) );
  AOI22_X1 U343 ( .A1(B[27]), .A2(n1413), .B1(A[27]), .B2(n1407), .ZN(n187) );
  AOI22_X1 U344 ( .A1(D[27]), .A2(n1425), .B1(C[27]), .B2(n1419), .ZN(n188) );
  AOI22_X1 U345 ( .A1(H[27]), .A2(n1449), .B1(G[27]), .B2(n1443), .ZN(n190) );
  NAND4_X1 U346 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U347 ( .A1(B[35]), .A2(n1414), .B1(A[35]), .B2(n1408), .ZN(n151) );
  AOI22_X1 U348 ( .A1(D[35]), .A2(n1426), .B1(C[35]), .B2(n1420), .ZN(n152) );
  AOI22_X1 U349 ( .A1(H[35]), .A2(n1450), .B1(G[35]), .B2(n1444), .ZN(n154) );
  AOI22_X1 U350 ( .A1(F[37]), .A2(n1438), .B1(E[37]), .B2(n1432), .ZN(n145) );
  AOI22_X1 U351 ( .A1(F[31]), .A2(n1438), .B1(E[31]), .B2(n1432), .ZN(n169) );
  NAND4_X1 U352 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U353 ( .A1(B[2]), .A2(n1413), .B1(A[2]), .B2(n1407), .ZN(n175) );
  AOI22_X1 U354 ( .A1(D[2]), .A2(n1425), .B1(C[2]), .B2(n1419), .ZN(n176) );
  AOI22_X1 U355 ( .A1(F[2]), .A2(n1437), .B1(E[2]), .B2(n1431), .ZN(n177) );
  NAND4_X1 U356 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U357 ( .A1(B[0]), .A2(n1412), .B1(A[0]), .B2(n1406), .ZN(n263) );
  AOI22_X1 U358 ( .A1(D[0]), .A2(n1424), .B1(C[0]), .B2(n1418), .ZN(n264) );
  AOI22_X1 U359 ( .A1(F[0]), .A2(n1436), .B1(E[0]), .B2(n1430), .ZN(n265) );
  AOI22_X1 U360 ( .A1(H[3]), .A2(n1450), .B1(G[3]), .B2(n1444), .ZN(n134) );
  AOI22_X1 U361 ( .A1(H[2]), .A2(n1449), .B1(G[2]), .B2(n1443), .ZN(n178) );
  AOI22_X1 U362 ( .A1(H[1]), .A2(n1448), .B1(G[1]), .B2(n1442), .ZN(n222) );
  NAND4_X1 U363 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U364 ( .A1(B[3]), .A2(n1414), .B1(A[3]), .B2(n1408), .ZN(n131) );
  AOI22_X1 U365 ( .A1(D[3]), .A2(n1426), .B1(C[3]), .B2(n1420), .ZN(n132) );
  AOI22_X1 U366 ( .A1(F[3]), .A2(n1438), .B1(E[3]), .B2(n1432), .ZN(n133) );
  NAND4_X1 U367 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U368 ( .A1(B[1]), .A2(n1412), .B1(A[1]), .B2(n1406), .ZN(n219) );
  AOI22_X1 U369 ( .A1(D[1]), .A2(n1424), .B1(C[1]), .B2(n1418), .ZN(n220) );
  AOI22_X1 U370 ( .A1(F[1]), .A2(n1436), .B1(E[1]), .B2(n1430), .ZN(n221) );
  AOI22_X1 U371 ( .A1(H[0]), .A2(n1448), .B1(G[0]), .B2(n1442), .ZN(n266) );
  CLKBUF_X1 U372 ( .A(n14), .Z(n1411) );
  CLKBUF_X1 U373 ( .A(n13), .Z(n1417) );
  CLKBUF_X1 U374 ( .A(n12), .Z(n1423) );
  CLKBUF_X1 U375 ( .A(n11), .Z(n1429) );
  CLKBUF_X1 U376 ( .A(n10), .Z(n1435) );
  CLKBUF_X1 U377 ( .A(n9), .Z(n1441) );
  CLKBUF_X1 U378 ( .A(n8), .Z(n1447) );
  CLKBUF_X1 U379 ( .A(n7), .Z(n1453) );
endmodule


module MUX81_GENERIC_NBIT64_13 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444;

  BUF_X1 U1 ( .A(n13), .Z(n1401) );
  BUF_X1 U2 ( .A(n13), .Z(n1402) );
  BUF_X1 U3 ( .A(n13), .Z(n1403) );
  BUF_X1 U4 ( .A(n12), .Z(n1408) );
  BUF_X1 U5 ( .A(n12), .Z(n1407) );
  BUF_X1 U6 ( .A(n12), .Z(n1409) );
  BUF_X1 U7 ( .A(n10), .Z(n1419) );
  BUF_X1 U8 ( .A(n8), .Z(n1431) );
  BUF_X1 U9 ( .A(n8), .Z(n1432) );
  BUF_X1 U10 ( .A(n8), .Z(n1433) );
  BUF_X1 U11 ( .A(n10), .Z(n1420) );
  BUF_X1 U12 ( .A(n10), .Z(n1421) );
  BUF_X1 U13 ( .A(n13), .Z(n1404) );
  BUF_X1 U14 ( .A(n12), .Z(n1410) );
  BUF_X1 U15 ( .A(n12), .Z(n1411) );
  BUF_X1 U16 ( .A(n8), .Z(n1434) );
  BUF_X1 U17 ( .A(n10), .Z(n1422) );
  BUF_X1 U18 ( .A(n10), .Z(n1423) );
  BUF_X1 U19 ( .A(n13), .Z(n1405) );
  BUF_X1 U20 ( .A(n8), .Z(n1435) );
  BUF_X1 U21 ( .A(n11), .Z(n1416) );
  BUF_X1 U22 ( .A(n11), .Z(n1414) );
  BUF_X1 U23 ( .A(n11), .Z(n1415) );
  BUF_X1 U24 ( .A(n11), .Z(n1413) );
  BUF_X1 U25 ( .A(n11), .Z(n1417) );
  BUF_X1 U26 ( .A(n7), .Z(n1437) );
  BUF_X1 U27 ( .A(n7), .Z(n1438) );
  BUF_X1 U28 ( .A(n7), .Z(n1439) );
  BUF_X1 U29 ( .A(n7), .Z(n1440) );
  BUF_X1 U30 ( .A(n9), .Z(n1428) );
  BUF_X1 U31 ( .A(n7), .Z(n1441) );
  BUF_X1 U32 ( .A(n9), .Z(n1426) );
  BUF_X1 U33 ( .A(n9), .Z(n1427) );
  BUF_X1 U34 ( .A(n9), .Z(n1425) );
  BUF_X1 U35 ( .A(n9), .Z(n1429) );
  BUF_X1 U36 ( .A(n14), .Z(n1398) );
  BUF_X1 U37 ( .A(n14), .Z(n1396) );
  BUF_X1 U38 ( .A(n14), .Z(n1397) );
  BUF_X1 U39 ( .A(n14), .Z(n1395) );
  BUF_X1 U40 ( .A(n14), .Z(n1399) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1443), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1444), .ZN(n13) );
  AND3_X1 U43 ( .A1(n1444), .A2(n1443), .A3(SEL[2]), .ZN(n10) );
  AND3_X1 U44 ( .A1(SEL[1]), .A2(n1444), .A3(SEL[2]), .ZN(n8) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1443) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1444) );
  NOR3_X1 U47 ( .A1(n1444), .A2(SEL[2]), .A3(n1443), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1443), .A3(SEL[2]), .ZN(n9) );
  AOI22_X1 U51 ( .A1(H[22]), .A2(n1438), .B1(G[22]), .B2(n1432), .ZN(n210) );
  AOI22_X1 U52 ( .A1(H[42]), .A2(n1440), .B1(G[42]), .B2(n1434), .ZN(n122) );
  NAND4_X1 U53 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U54 ( .A1(B[14]), .A2(n1401), .B1(A[14]), .B2(n1395), .ZN(n243) );
  AOI22_X1 U55 ( .A1(H[14]), .A2(n1437), .B1(G[14]), .B2(n1431), .ZN(n246) );
  AOI22_X1 U56 ( .A1(D[14]), .A2(n1413), .B1(C[14]), .B2(n1407), .ZN(n244) );
  NAND4_X1 U57 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U58 ( .A1(H[10]), .A2(n1437), .B1(G[10]), .B2(n1431), .ZN(n262) );
  AOI22_X1 U59 ( .A1(B[10]), .A2(n1401), .B1(A[10]), .B2(n1395), .ZN(n259) );
  AOI22_X1 U60 ( .A1(D[10]), .A2(n1413), .B1(C[10]), .B2(n1407), .ZN(n260) );
  NAND4_X1 U61 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U62 ( .A1(H[8]), .A2(n1442), .B1(G[8]), .B2(n1436), .ZN(n18) );
  AOI22_X1 U63 ( .A1(B[8]), .A2(n1406), .B1(A[8]), .B2(n1400), .ZN(n15) );
  AOI22_X1 U64 ( .A1(D[8]), .A2(n1418), .B1(C[8]), .B2(n1412), .ZN(n16) );
  NAND4_X1 U65 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U66 ( .A1(B[17]), .A2(n1401), .B1(A[17]), .B2(n1395), .ZN(n231) );
  AOI22_X1 U67 ( .A1(D[17]), .A2(n1413), .B1(C[17]), .B2(n1407), .ZN(n232) );
  AOI22_X1 U68 ( .A1(F[17]), .A2(n1425), .B1(E[17]), .B2(n1419), .ZN(n233) );
  AOI22_X1 U69 ( .A1(H[37]), .A2(n1439), .B1(G[37]), .B2(n1433), .ZN(n146) );
  AOI22_X1 U70 ( .A1(H[36]), .A2(n1439), .B1(G[36]), .B2(n1433), .ZN(n150) );
  AOI22_X1 U71 ( .A1(H[40]), .A2(n1439), .B1(G[40]), .B2(n1433), .ZN(n130) );
  AOI22_X1 U72 ( .A1(H[33]), .A2(n1439), .B1(G[33]), .B2(n1433), .ZN(n162) );
  AOI22_X1 U73 ( .A1(H[38]), .A2(n1439), .B1(G[38]), .B2(n1433), .ZN(n142) );
  AOI22_X1 U74 ( .A1(H[35]), .A2(n1439), .B1(G[35]), .B2(n1433), .ZN(n154) );
  AOI22_X1 U75 ( .A1(H[34]), .A2(n1439), .B1(G[34]), .B2(n1433), .ZN(n158) );
  AOI22_X1 U76 ( .A1(H[48]), .A2(n1440), .B1(G[48]), .B2(n1434), .ZN(n98) );
  AOI22_X1 U77 ( .A1(H[54]), .A2(n1441), .B1(G[54]), .B2(n1435), .ZN(n70) );
  AOI22_X1 U78 ( .A1(H[56]), .A2(n1441), .B1(G[56]), .B2(n1435), .ZN(n62) );
  AOI22_X1 U79 ( .A1(H[44]), .A2(n1440), .B1(G[44]), .B2(n1434), .ZN(n114) );
  AOI22_X1 U80 ( .A1(H[45]), .A2(n1440), .B1(G[45]), .B2(n1434), .ZN(n110) );
  AOI22_X1 U81 ( .A1(H[46]), .A2(n1440), .B1(G[46]), .B2(n1434), .ZN(n106) );
  AOI22_X1 U82 ( .A1(H[52]), .A2(n1440), .B1(G[52]), .B2(n1434), .ZN(n78) );
  AOI22_X1 U83 ( .A1(H[32]), .A2(n1439), .B1(G[32]), .B2(n1433), .ZN(n166) );
  AOI22_X1 U84 ( .A1(H[29]), .A2(n1438), .B1(G[29]), .B2(n1432), .ZN(n182) );
  AOI22_X1 U85 ( .A1(H[39]), .A2(n1439), .B1(G[39]), .B2(n1433), .ZN(n138) );
  AOI22_X1 U86 ( .A1(H[49]), .A2(n1440), .B1(G[49]), .B2(n1434), .ZN(n94) );
  AOI22_X1 U87 ( .A1(H[47]), .A2(n1440), .B1(G[47]), .B2(n1434), .ZN(n102) );
  AOI22_X1 U88 ( .A1(H[30]), .A2(n1438), .B1(G[30]), .B2(n1432), .ZN(n174) );
  AOI22_X1 U89 ( .A1(H[50]), .A2(n1440), .B1(G[50]), .B2(n1434), .ZN(n86) );
  AOI22_X1 U90 ( .A1(H[31]), .A2(n1439), .B1(G[31]), .B2(n1433), .ZN(n170) );
  AOI22_X1 U91 ( .A1(H[57]), .A2(n1441), .B1(G[57]), .B2(n1435), .ZN(n58) );
  AOI22_X1 U92 ( .A1(H[55]), .A2(n1441), .B1(G[55]), .B2(n1435), .ZN(n66) );
  AOI22_X1 U93 ( .A1(H[53]), .A2(n1441), .B1(G[53]), .B2(n1435), .ZN(n74) );
  AOI22_X1 U94 ( .A1(H[51]), .A2(n1440), .B1(G[51]), .B2(n1434), .ZN(n82) );
  AOI22_X1 U95 ( .A1(H[58]), .A2(n1441), .B1(G[58]), .B2(n1435), .ZN(n54) );
  AOI22_X1 U96 ( .A1(H[28]), .A2(n1438), .B1(G[28]), .B2(n1432), .ZN(n186) );
  AOI22_X1 U97 ( .A1(H[60]), .A2(n1441), .B1(G[60]), .B2(n1435), .ZN(n42) );
  AOI22_X1 U98 ( .A1(H[27]), .A2(n1438), .B1(G[27]), .B2(n1432), .ZN(n190) );
  AOI22_X1 U99 ( .A1(H[26]), .A2(n1438), .B1(G[26]), .B2(n1432), .ZN(n194) );
  AOI22_X1 U100 ( .A1(H[24]), .A2(n1438), .B1(G[24]), .B2(n1432), .ZN(n202) );
  AOI22_X1 U101 ( .A1(H[25]), .A2(n1438), .B1(G[25]), .B2(n1432), .ZN(n198) );
  AOI22_X1 U102 ( .A1(H[21]), .A2(n1438), .B1(G[21]), .B2(n1432), .ZN(n214) );
  AOI22_X1 U103 ( .A1(H[59]), .A2(n1441), .B1(G[59]), .B2(n1435), .ZN(n50) );
  AOI22_X1 U104 ( .A1(H[20]), .A2(n1438), .B1(G[20]), .B2(n1432), .ZN(n218) );
  AOI22_X1 U105 ( .A1(H[23]), .A2(n1438), .B1(G[23]), .B2(n1432), .ZN(n206) );
  AOI22_X1 U106 ( .A1(H[17]), .A2(n1437), .B1(G[17]), .B2(n1431), .ZN(n234) );
  AOI22_X1 U107 ( .A1(H[16]), .A2(n1437), .B1(G[16]), .B2(n1431), .ZN(n238) );
  AOI22_X1 U108 ( .A1(H[18]), .A2(n1437), .B1(G[18]), .B2(n1431), .ZN(n230) );
  AOI22_X1 U109 ( .A1(H[19]), .A2(n1437), .B1(G[19]), .B2(n1431), .ZN(n226) );
  AOI22_X1 U110 ( .A1(H[61]), .A2(n1441), .B1(G[61]), .B2(n1435), .ZN(n38) );
  AOI22_X1 U111 ( .A1(H[62]), .A2(n1441), .B1(G[62]), .B2(n1435), .ZN(n34) );
  AOI22_X1 U112 ( .A1(H[63]), .A2(n1441), .B1(G[63]), .B2(n1435), .ZN(n30) );
  NAND4_X1 U113 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U114 ( .A1(B[21]), .A2(n1402), .B1(A[21]), .B2(n1396), .ZN(n211) );
  AOI22_X1 U115 ( .A1(D[21]), .A2(n1414), .B1(C[21]), .B2(n1408), .ZN(n212) );
  AOI22_X1 U116 ( .A1(F[21]), .A2(n1426), .B1(E[21]), .B2(n1420), .ZN(n213) );
  AOI22_X1 U117 ( .A1(F[10]), .A2(n1425), .B1(E[10]), .B2(n1419), .ZN(n261) );
  AOI22_X1 U118 ( .A1(F[15]), .A2(n1425), .B1(E[15]), .B2(n1419), .ZN(n241) );
  AOI22_X1 U119 ( .A1(F[13]), .A2(n1425), .B1(E[13]), .B2(n1419), .ZN(n249) );
  AOI22_X1 U120 ( .A1(F[14]), .A2(n1425), .B1(E[14]), .B2(n1419), .ZN(n245) );
  AOI22_X1 U121 ( .A1(F[8]), .A2(n1430), .B1(E[8]), .B2(n1424), .ZN(n17) );
  AOI22_X1 U122 ( .A1(F[6]), .A2(n1430), .B1(E[6]), .B2(n1424), .ZN(n25) );
  NAND4_X1 U123 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U124 ( .A1(H[11]), .A2(n1437), .B1(G[11]), .B2(n1431), .ZN(n258) );
  AOI22_X1 U125 ( .A1(B[11]), .A2(n1401), .B1(A[11]), .B2(n1395), .ZN(n255) );
  AOI22_X1 U126 ( .A1(F[11]), .A2(n1425), .B1(E[11]), .B2(n1419), .ZN(n257) );
  AOI22_X1 U127 ( .A1(D[11]), .A2(n1413), .B1(C[11]), .B2(n1407), .ZN(n256) );
  AOI22_X1 U128 ( .A1(D[12]), .A2(n1413), .B1(C[12]), .B2(n1407), .ZN(n252) );
  AOI22_X1 U129 ( .A1(D[9]), .A2(n1418), .B1(C[9]), .B2(n1412), .ZN(n4) );
  AOI22_X1 U130 ( .A1(D[7]), .A2(n1418), .B1(C[7]), .B2(n1412), .ZN(n20) );
  NAND4_X1 U131 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U132 ( .A1(H[9]), .A2(n1442), .B1(G[9]), .B2(n1436), .ZN(n6) );
  AOI22_X1 U133 ( .A1(B[9]), .A2(n1406), .B1(A[9]), .B2(n1400), .ZN(n3) );
  AOI22_X1 U134 ( .A1(F[9]), .A2(n1430), .B1(E[9]), .B2(n1424), .ZN(n5) );
  NAND4_X1 U135 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U136 ( .A1(B[27]), .A2(n1402), .B1(A[27]), .B2(n1396), .ZN(n187) );
  AOI22_X1 U137 ( .A1(D[27]), .A2(n1414), .B1(C[27]), .B2(n1408), .ZN(n188) );
  AOI22_X1 U138 ( .A1(F[27]), .A2(n1426), .B1(E[27]), .B2(n1420), .ZN(n189) );
  NAND4_X1 U139 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U140 ( .A1(B[26]), .A2(n1402), .B1(A[26]), .B2(n1396), .ZN(n191) );
  AOI22_X1 U141 ( .A1(D[26]), .A2(n1414), .B1(C[26]), .B2(n1408), .ZN(n192) );
  AOI22_X1 U142 ( .A1(F[26]), .A2(n1426), .B1(E[26]), .B2(n1420), .ZN(n193) );
  NAND4_X1 U143 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U144 ( .A1(B[15]), .A2(n1401), .B1(A[15]), .B2(n1395), .ZN(n239) );
  AOI22_X1 U145 ( .A1(H[15]), .A2(n1437), .B1(G[15]), .B2(n1431), .ZN(n242) );
  AOI22_X1 U146 ( .A1(D[15]), .A2(n1413), .B1(C[15]), .B2(n1407), .ZN(n240) );
  NAND4_X1 U147 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U148 ( .A1(B[23]), .A2(n1402), .B1(A[23]), .B2(n1396), .ZN(n203) );
  AOI22_X1 U149 ( .A1(D[23]), .A2(n1414), .B1(C[23]), .B2(n1408), .ZN(n204) );
  AOI22_X1 U150 ( .A1(F[23]), .A2(n1426), .B1(E[23]), .B2(n1420), .ZN(n205) );
  NAND4_X1 U151 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U152 ( .A1(B[18]), .A2(n1401), .B1(A[18]), .B2(n1395), .ZN(n227) );
  AOI22_X1 U153 ( .A1(D[18]), .A2(n1413), .B1(C[18]), .B2(n1407), .ZN(n228) );
  AOI22_X1 U154 ( .A1(F[18]), .A2(n1425), .B1(E[18]), .B2(n1419), .ZN(n229) );
  NAND4_X1 U155 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U156 ( .A1(B[19]), .A2(n1401), .B1(A[19]), .B2(n1395), .ZN(n223) );
  AOI22_X1 U157 ( .A1(D[19]), .A2(n1413), .B1(C[19]), .B2(n1407), .ZN(n224) );
  AOI22_X1 U158 ( .A1(F[19]), .A2(n1425), .B1(E[19]), .B2(n1419), .ZN(n225) );
  NAND4_X1 U159 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U160 ( .A1(B[16]), .A2(n1401), .B1(A[16]), .B2(n1395), .ZN(n235) );
  AOI22_X1 U161 ( .A1(D[16]), .A2(n1413), .B1(C[16]), .B2(n1407), .ZN(n236) );
  AOI22_X1 U162 ( .A1(F[16]), .A2(n1425), .B1(E[16]), .B2(n1419), .ZN(n237) );
  NAND4_X1 U163 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U164 ( .A1(B[33]), .A2(n1403), .B1(A[33]), .B2(n1397), .ZN(n159) );
  AOI22_X1 U165 ( .A1(D[33]), .A2(n1415), .B1(C[33]), .B2(n1409), .ZN(n160) );
  AOI22_X1 U166 ( .A1(F[33]), .A2(n1427), .B1(E[33]), .B2(n1421), .ZN(n161) );
  NAND4_X1 U167 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U168 ( .A1(B[37]), .A2(n1403), .B1(A[37]), .B2(n1397), .ZN(n143) );
  AOI22_X1 U169 ( .A1(D[37]), .A2(n1415), .B1(C[37]), .B2(n1409), .ZN(n144) );
  AOI22_X1 U170 ( .A1(F[37]), .A2(n1427), .B1(E[37]), .B2(n1421), .ZN(n145) );
  NAND4_X1 U171 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U172 ( .A1(B[34]), .A2(n1403), .B1(A[34]), .B2(n1397), .ZN(n155) );
  AOI22_X1 U173 ( .A1(D[34]), .A2(n1415), .B1(C[34]), .B2(n1409), .ZN(n156) );
  AOI22_X1 U174 ( .A1(F[34]), .A2(n1427), .B1(E[34]), .B2(n1421), .ZN(n157) );
  NAND4_X1 U175 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U176 ( .A1(B[32]), .A2(n1403), .B1(A[32]), .B2(n1397), .ZN(n163) );
  AOI22_X1 U177 ( .A1(D[32]), .A2(n1415), .B1(C[32]), .B2(n1409), .ZN(n164) );
  AOI22_X1 U178 ( .A1(F[32]), .A2(n1427), .B1(E[32]), .B2(n1421), .ZN(n165) );
  NAND4_X1 U179 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U180 ( .A1(B[29]), .A2(n1402), .B1(A[29]), .B2(n1396), .ZN(n179) );
  AOI22_X1 U181 ( .A1(D[29]), .A2(n1414), .B1(C[29]), .B2(n1408), .ZN(n180) );
  AOI22_X1 U182 ( .A1(F[29]), .A2(n1426), .B1(E[29]), .B2(n1420), .ZN(n181) );
  NAND4_X1 U183 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U184 ( .A1(B[36]), .A2(n1403), .B1(A[36]), .B2(n1397), .ZN(n147) );
  AOI22_X1 U185 ( .A1(D[36]), .A2(n1415), .B1(C[36]), .B2(n1409), .ZN(n148) );
  AOI22_X1 U186 ( .A1(F[36]), .A2(n1427), .B1(E[36]), .B2(n1421), .ZN(n149) );
  NAND4_X1 U187 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U188 ( .A1(B[40]), .A2(n1403), .B1(A[40]), .B2(n1397), .ZN(n127) );
  AOI22_X1 U189 ( .A1(D[40]), .A2(n1415), .B1(C[40]), .B2(n1409), .ZN(n128) );
  AOI22_X1 U190 ( .A1(F[40]), .A2(n1427), .B1(E[40]), .B2(n1421), .ZN(n129) );
  NAND4_X1 U191 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U192 ( .A1(B[28]), .A2(n1402), .B1(A[28]), .B2(n1396), .ZN(n183) );
  AOI22_X1 U193 ( .A1(D[28]), .A2(n1414), .B1(C[28]), .B2(n1408), .ZN(n184) );
  AOI22_X1 U194 ( .A1(F[28]), .A2(n1426), .B1(E[28]), .B2(n1420), .ZN(n185) );
  NAND4_X1 U195 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U196 ( .A1(B[38]), .A2(n1403), .B1(A[38]), .B2(n1397), .ZN(n139) );
  AOI22_X1 U197 ( .A1(D[38]), .A2(n1415), .B1(C[38]), .B2(n1409), .ZN(n140) );
  AOI22_X1 U198 ( .A1(F[38]), .A2(n1427), .B1(E[38]), .B2(n1421), .ZN(n141) );
  NAND4_X1 U199 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U200 ( .A1(B[41]), .A2(n1403), .B1(A[41]), .B2(n1397), .ZN(n123) );
  AOI22_X1 U201 ( .A1(D[41]), .A2(n1415), .B1(C[41]), .B2(n1409), .ZN(n124) );
  AOI22_X1 U202 ( .A1(F[41]), .A2(n1427), .B1(E[41]), .B2(n1421), .ZN(n125) );
  NAND4_X1 U203 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U204 ( .A1(B[24]), .A2(n1402), .B1(A[24]), .B2(n1396), .ZN(n199) );
  AOI22_X1 U205 ( .A1(D[24]), .A2(n1414), .B1(C[24]), .B2(n1408), .ZN(n200) );
  AOI22_X1 U206 ( .A1(F[24]), .A2(n1426), .B1(E[24]), .B2(n1420), .ZN(n201) );
  NAND4_X1 U207 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U208 ( .A1(B[48]), .A2(n1404), .B1(A[48]), .B2(n1398), .ZN(n95) );
  AOI22_X1 U209 ( .A1(D[48]), .A2(n1416), .B1(C[48]), .B2(n1410), .ZN(n96) );
  AOI22_X1 U210 ( .A1(F[48]), .A2(n1428), .B1(E[48]), .B2(n1422), .ZN(n97) );
  NAND4_X1 U211 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U212 ( .A1(B[54]), .A2(n1405), .B1(A[54]), .B2(n1399), .ZN(n67) );
  AOI22_X1 U213 ( .A1(D[54]), .A2(n1417), .B1(C[54]), .B2(n1411), .ZN(n68) );
  AOI22_X1 U214 ( .A1(F[54]), .A2(n1429), .B1(E[54]), .B2(n1423), .ZN(n69) );
  NAND4_X1 U215 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U216 ( .A1(B[56]), .A2(n1405), .B1(A[56]), .B2(n1399), .ZN(n59) );
  AOI22_X1 U217 ( .A1(D[56]), .A2(n1417), .B1(C[56]), .B2(n1411), .ZN(n60) );
  AOI22_X1 U218 ( .A1(F[56]), .A2(n1429), .B1(E[56]), .B2(n1423), .ZN(n61) );
  NAND4_X1 U219 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U220 ( .A1(B[42]), .A2(n1404), .B1(A[42]), .B2(n1398), .ZN(n119) );
  AOI22_X1 U221 ( .A1(D[42]), .A2(n1416), .B1(C[42]), .B2(n1410), .ZN(n120) );
  AOI22_X1 U222 ( .A1(F[42]), .A2(n1428), .B1(E[42]), .B2(n1422), .ZN(n121) );
  NAND4_X1 U223 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U224 ( .A1(B[44]), .A2(n1404), .B1(A[44]), .B2(n1398), .ZN(n111) );
  AOI22_X1 U225 ( .A1(D[44]), .A2(n1416), .B1(C[44]), .B2(n1410), .ZN(n112) );
  AOI22_X1 U226 ( .A1(F[44]), .A2(n1428), .B1(E[44]), .B2(n1422), .ZN(n113) );
  NAND4_X1 U227 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U228 ( .A1(B[45]), .A2(n1404), .B1(A[45]), .B2(n1398), .ZN(n107) );
  AOI22_X1 U229 ( .A1(D[45]), .A2(n1416), .B1(C[45]), .B2(n1410), .ZN(n108) );
  AOI22_X1 U230 ( .A1(F[45]), .A2(n1428), .B1(E[45]), .B2(n1422), .ZN(n109) );
  NAND4_X1 U231 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U232 ( .A1(B[46]), .A2(n1404), .B1(A[46]), .B2(n1398), .ZN(n103) );
  AOI22_X1 U233 ( .A1(D[46]), .A2(n1416), .B1(C[46]), .B2(n1410), .ZN(n104) );
  AOI22_X1 U234 ( .A1(F[46]), .A2(n1428), .B1(E[46]), .B2(n1422), .ZN(n105) );
  NAND4_X1 U235 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U236 ( .A1(B[20]), .A2(n1402), .B1(A[20]), .B2(n1396), .ZN(n215) );
  AOI22_X1 U237 ( .A1(D[20]), .A2(n1414), .B1(C[20]), .B2(n1408), .ZN(n216) );
  AOI22_X1 U238 ( .A1(F[20]), .A2(n1426), .B1(E[20]), .B2(n1420), .ZN(n217) );
  NAND4_X1 U239 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U240 ( .A1(B[52]), .A2(n1404), .B1(A[52]), .B2(n1398), .ZN(n75) );
  AOI22_X1 U241 ( .A1(D[52]), .A2(n1416), .B1(C[52]), .B2(n1410), .ZN(n76) );
  AOI22_X1 U242 ( .A1(F[52]), .A2(n1428), .B1(E[52]), .B2(n1422), .ZN(n77) );
  NAND4_X1 U243 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U244 ( .A1(B[49]), .A2(n1404), .B1(A[49]), .B2(n1398), .ZN(n91) );
  AOI22_X1 U245 ( .A1(D[49]), .A2(n1416), .B1(C[49]), .B2(n1410), .ZN(n92) );
  AOI22_X1 U246 ( .A1(F[49]), .A2(n1428), .B1(E[49]), .B2(n1422), .ZN(n93) );
  NAND4_X1 U247 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U248 ( .A1(H[12]), .A2(n1437), .B1(G[12]), .B2(n1431), .ZN(n254) );
  AOI22_X1 U249 ( .A1(B[12]), .A2(n1401), .B1(A[12]), .B2(n1395), .ZN(n251) );
  AOI22_X1 U250 ( .A1(F[12]), .A2(n1425), .B1(E[12]), .B2(n1419), .ZN(n253) );
  NAND4_X1 U251 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U252 ( .A1(B[50]), .A2(n1404), .B1(A[50]), .B2(n1398), .ZN(n83) );
  AOI22_X1 U253 ( .A1(D[50]), .A2(n1416), .B1(C[50]), .B2(n1410), .ZN(n84) );
  AOI22_X1 U254 ( .A1(F[50]), .A2(n1428), .B1(E[50]), .B2(n1422), .ZN(n85) );
  NAND4_X1 U255 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U256 ( .A1(B[57]), .A2(n1405), .B1(A[57]), .B2(n1399), .ZN(n55) );
  AOI22_X1 U257 ( .A1(D[57]), .A2(n1417), .B1(C[57]), .B2(n1411), .ZN(n56) );
  AOI22_X1 U258 ( .A1(F[57]), .A2(n1429), .B1(E[57]), .B2(n1423), .ZN(n57) );
  NAND4_X1 U259 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U260 ( .A1(B[53]), .A2(n1405), .B1(A[53]), .B2(n1399), .ZN(n71) );
  AOI22_X1 U261 ( .A1(D[53]), .A2(n1417), .B1(C[53]), .B2(n1411), .ZN(n72) );
  AOI22_X1 U262 ( .A1(F[53]), .A2(n1429), .B1(E[53]), .B2(n1423), .ZN(n73) );
  NAND4_X1 U263 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U264 ( .A1(B[58]), .A2(n1405), .B1(A[58]), .B2(n1399), .ZN(n51) );
  AOI22_X1 U265 ( .A1(D[58]), .A2(n1417), .B1(C[58]), .B2(n1411), .ZN(n52) );
  AOI22_X1 U266 ( .A1(F[58]), .A2(n1429), .B1(E[58]), .B2(n1423), .ZN(n53) );
  NAND4_X1 U267 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U268 ( .A1(B[60]), .A2(n1405), .B1(A[60]), .B2(n1399), .ZN(n39) );
  AOI22_X1 U269 ( .A1(D[60]), .A2(n1417), .B1(C[60]), .B2(n1411), .ZN(n40) );
  AOI22_X1 U270 ( .A1(F[60]), .A2(n1429), .B1(E[60]), .B2(n1423), .ZN(n41) );
  NAND4_X1 U271 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U272 ( .A1(B[61]), .A2(n1405), .B1(A[61]), .B2(n1399), .ZN(n35) );
  AOI22_X1 U273 ( .A1(D[61]), .A2(n1417), .B1(C[61]), .B2(n1411), .ZN(n36) );
  AOI22_X1 U274 ( .A1(F[61]), .A2(n1429), .B1(E[61]), .B2(n1423), .ZN(n37) );
  NAND4_X1 U275 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U276 ( .A1(B[62]), .A2(n1405), .B1(A[62]), .B2(n1399), .ZN(n31) );
  AOI22_X1 U277 ( .A1(D[62]), .A2(n1417), .B1(C[62]), .B2(n1411), .ZN(n32) );
  AOI22_X1 U278 ( .A1(F[62]), .A2(n1429), .B1(E[62]), .B2(n1423), .ZN(n33) );
  NAND4_X1 U279 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U280 ( .A1(B[63]), .A2(n1405), .B1(A[63]), .B2(n1399), .ZN(n27) );
  AOI22_X1 U281 ( .A1(D[63]), .A2(n1417), .B1(C[63]), .B2(n1411), .ZN(n28) );
  AOI22_X1 U282 ( .A1(F[63]), .A2(n1429), .B1(E[63]), .B2(n1423), .ZN(n29) );
  NAND4_X1 U283 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U284 ( .A1(D[6]), .A2(n1418), .B1(C[6]), .B2(n1412), .ZN(n24) );
  AOI22_X1 U285 ( .A1(H[6]), .A2(n1442), .B1(G[6]), .B2(n1436), .ZN(n26) );
  AOI22_X1 U286 ( .A1(B[6]), .A2(n1406), .B1(A[6]), .B2(n1400), .ZN(n23) );
  NAND4_X1 U287 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U288 ( .A1(H[13]), .A2(n1437), .B1(G[13]), .B2(n1431), .ZN(n250) );
  AOI22_X1 U289 ( .A1(B[13]), .A2(n1401), .B1(A[13]), .B2(n1395), .ZN(n247) );
  AOI22_X1 U290 ( .A1(D[13]), .A2(n1413), .B1(C[13]), .B2(n1407), .ZN(n248) );
  NAND4_X1 U291 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U292 ( .A1(H[7]), .A2(n1442), .B1(G[7]), .B2(n1436), .ZN(n22) );
  AOI22_X1 U293 ( .A1(B[7]), .A2(n1406), .B1(A[7]), .B2(n1400), .ZN(n19) );
  AOI22_X1 U294 ( .A1(F[7]), .A2(n1430), .B1(E[7]), .B2(n1424), .ZN(n21) );
  AOI22_X1 U295 ( .A1(H[43]), .A2(n1440), .B1(G[43]), .B2(n1434), .ZN(n118) );
  NAND4_X1 U296 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U297 ( .A1(B[47]), .A2(n1404), .B1(A[47]), .B2(n1398), .ZN(n99) );
  AOI22_X1 U298 ( .A1(D[47]), .A2(n1416), .B1(C[47]), .B2(n1410), .ZN(n100) );
  AOI22_X1 U299 ( .A1(F[47]), .A2(n1428), .B1(E[47]), .B2(n1422), .ZN(n101) );
  AOI22_X1 U300 ( .A1(H[41]), .A2(n1439), .B1(G[41]), .B2(n1433), .ZN(n126) );
  NAND4_X1 U301 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U302 ( .A1(B[31]), .A2(n1403), .B1(A[31]), .B2(n1397), .ZN(n167) );
  AOI22_X1 U303 ( .A1(D[31]), .A2(n1415), .B1(C[31]), .B2(n1409), .ZN(n168) );
  AOI22_X1 U304 ( .A1(F[31]), .A2(n1427), .B1(E[31]), .B2(n1421), .ZN(n169) );
  NAND4_X1 U305 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U306 ( .A1(B[55]), .A2(n1405), .B1(A[55]), .B2(n1399), .ZN(n63) );
  AOI22_X1 U307 ( .A1(D[55]), .A2(n1417), .B1(C[55]), .B2(n1411), .ZN(n64) );
  AOI22_X1 U308 ( .A1(F[55]), .A2(n1429), .B1(E[55]), .B2(n1423), .ZN(n65) );
  NAND4_X1 U309 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U310 ( .A1(B[59]), .A2(n1405), .B1(A[59]), .B2(n1399), .ZN(n47) );
  AOI22_X1 U311 ( .A1(D[59]), .A2(n1417), .B1(C[59]), .B2(n1411), .ZN(n48) );
  AOI22_X1 U312 ( .A1(F[59]), .A2(n1429), .B1(E[59]), .B2(n1423), .ZN(n49) );
  NAND4_X1 U313 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U314 ( .A1(B[35]), .A2(n1403), .B1(A[35]), .B2(n1397), .ZN(n151) );
  AOI22_X1 U315 ( .A1(D[35]), .A2(n1415), .B1(C[35]), .B2(n1409), .ZN(n152) );
  AOI22_X1 U316 ( .A1(F[35]), .A2(n1427), .B1(E[35]), .B2(n1421), .ZN(n153) );
  NAND4_X1 U317 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U318 ( .A1(B[22]), .A2(n1402), .B1(A[22]), .B2(n1396), .ZN(n207) );
  AOI22_X1 U319 ( .A1(D[22]), .A2(n1414), .B1(C[22]), .B2(n1408), .ZN(n208) );
  AOI22_X1 U320 ( .A1(F[22]), .A2(n1426), .B1(E[22]), .B2(n1420), .ZN(n209) );
  NAND4_X1 U321 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U322 ( .A1(B[30]), .A2(n1402), .B1(A[30]), .B2(n1396), .ZN(n171) );
  AOI22_X1 U323 ( .A1(D[30]), .A2(n1414), .B1(C[30]), .B2(n1408), .ZN(n172) );
  AOI22_X1 U324 ( .A1(F[30]), .A2(n1426), .B1(E[30]), .B2(n1420), .ZN(n173) );
  NAND4_X1 U325 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U326 ( .A1(B[25]), .A2(n1402), .B1(A[25]), .B2(n1396), .ZN(n195) );
  AOI22_X1 U327 ( .A1(D[25]), .A2(n1414), .B1(C[25]), .B2(n1408), .ZN(n196) );
  AOI22_X1 U328 ( .A1(F[25]), .A2(n1426), .B1(E[25]), .B2(n1420), .ZN(n197) );
  NAND4_X1 U329 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U330 ( .A1(B[39]), .A2(n1403), .B1(A[39]), .B2(n1397), .ZN(n135) );
  AOI22_X1 U331 ( .A1(D[39]), .A2(n1415), .B1(C[39]), .B2(n1409), .ZN(n136) );
  AOI22_X1 U332 ( .A1(F[39]), .A2(n1427), .B1(E[39]), .B2(n1421), .ZN(n137) );
  NAND4_X1 U333 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U334 ( .A1(B[43]), .A2(n1404), .B1(A[43]), .B2(n1398), .ZN(n115) );
  AOI22_X1 U335 ( .A1(D[43]), .A2(n1416), .B1(C[43]), .B2(n1410), .ZN(n116) );
  AOI22_X1 U336 ( .A1(F[43]), .A2(n1428), .B1(E[43]), .B2(n1422), .ZN(n117) );
  NAND4_X1 U337 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U338 ( .A1(B[51]), .A2(n1404), .B1(A[51]), .B2(n1398), .ZN(n79) );
  AOI22_X1 U339 ( .A1(D[51]), .A2(n1416), .B1(C[51]), .B2(n1410), .ZN(n80) );
  AOI22_X1 U340 ( .A1(F[51]), .A2(n1428), .B1(E[51]), .B2(n1422), .ZN(n81) );
  NAND4_X1 U341 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U342 ( .A1(B[5]), .A2(n1405), .B1(A[5]), .B2(n1399), .ZN(n43) );
  AOI22_X1 U343 ( .A1(D[5]), .A2(n1417), .B1(C[5]), .B2(n1411), .ZN(n44) );
  AOI22_X1 U344 ( .A1(F[5]), .A2(n1429), .B1(E[5]), .B2(n1423), .ZN(n45) );
  NAND4_X1 U345 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U346 ( .A1(B[0]), .A2(n1401), .B1(A[0]), .B2(n1395), .ZN(n263) );
  AOI22_X1 U347 ( .A1(D[0]), .A2(n1413), .B1(C[0]), .B2(n1407), .ZN(n264) );
  AOI22_X1 U348 ( .A1(F[0]), .A2(n1425), .B1(E[0]), .B2(n1419), .ZN(n265) );
  AOI22_X1 U349 ( .A1(H[4]), .A2(n1440), .B1(G[4]), .B2(n1434), .ZN(n90) );
  AOI22_X1 U350 ( .A1(H[3]), .A2(n1439), .B1(G[3]), .B2(n1433), .ZN(n134) );
  AOI22_X1 U351 ( .A1(H[5]), .A2(n1441), .B1(G[5]), .B2(n1435), .ZN(n46) );
  AOI22_X1 U352 ( .A1(H[2]), .A2(n1438), .B1(G[2]), .B2(n1432), .ZN(n178) );
  AOI22_X1 U353 ( .A1(H[1]), .A2(n1437), .B1(G[1]), .B2(n1431), .ZN(n222) );
  NAND4_X1 U354 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U355 ( .A1(B[3]), .A2(n1403), .B1(A[3]), .B2(n1397), .ZN(n131) );
  AOI22_X1 U356 ( .A1(D[3]), .A2(n1415), .B1(C[3]), .B2(n1409), .ZN(n132) );
  AOI22_X1 U357 ( .A1(F[3]), .A2(n1427), .B1(E[3]), .B2(n1421), .ZN(n133) );
  NAND4_X1 U358 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U359 ( .A1(B[2]), .A2(n1402), .B1(A[2]), .B2(n1396), .ZN(n175) );
  AOI22_X1 U360 ( .A1(D[2]), .A2(n1414), .B1(C[2]), .B2(n1408), .ZN(n176) );
  AOI22_X1 U361 ( .A1(F[2]), .A2(n1426), .B1(E[2]), .B2(n1420), .ZN(n177) );
  NAND4_X1 U362 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U363 ( .A1(B[4]), .A2(n1404), .B1(A[4]), .B2(n1398), .ZN(n87) );
  AOI22_X1 U364 ( .A1(D[4]), .A2(n1416), .B1(C[4]), .B2(n1410), .ZN(n88) );
  AOI22_X1 U365 ( .A1(F[4]), .A2(n1428), .B1(E[4]), .B2(n1422), .ZN(n89) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1401), .B1(A[1]), .B2(n1395), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1413), .B1(C[1]), .B2(n1407), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1425), .B1(E[1]), .B2(n1419), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1437), .B1(G[0]), .B2(n1431), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1400) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1406) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1412) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1418) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1424) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1430) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1436) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1442) );
endmodule


module MUX81_GENERIC_NBIT64_12 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446;

  BUF_X1 U1 ( .A(n13), .Z(n1403) );
  BUF_X1 U2 ( .A(n13), .Z(n1404) );
  BUF_X1 U3 ( .A(n13), .Z(n1405) );
  BUF_X1 U4 ( .A(n12), .Z(n1409) );
  BUF_X1 U5 ( .A(n12), .Z(n1410) );
  BUF_X1 U6 ( .A(n12), .Z(n1411) );
  BUF_X1 U7 ( .A(n8), .Z(n1433) );
  BUF_X1 U8 ( .A(n10), .Z(n1421) );
  BUF_X1 U9 ( .A(n8), .Z(n1434) );
  BUF_X1 U10 ( .A(n8), .Z(n1435) );
  BUF_X1 U11 ( .A(n10), .Z(n1422) );
  BUF_X1 U12 ( .A(n10), .Z(n1423) );
  BUF_X1 U13 ( .A(n13), .Z(n1406) );
  BUF_X1 U14 ( .A(n12), .Z(n1412) );
  BUF_X1 U15 ( .A(n10), .Z(n1424) );
  BUF_X1 U16 ( .A(n8), .Z(n1436) );
  BUF_X1 U17 ( .A(n13), .Z(n1407) );
  BUF_X1 U18 ( .A(n12), .Z(n1413) );
  BUF_X1 U19 ( .A(n10), .Z(n1425) );
  BUF_X1 U20 ( .A(n8), .Z(n1437) );
  BUF_X1 U21 ( .A(n11), .Z(n1418) );
  BUF_X1 U22 ( .A(n11), .Z(n1416) );
  BUF_X1 U23 ( .A(n11), .Z(n1417) );
  BUF_X1 U24 ( .A(n11), .Z(n1415) );
  BUF_X1 U25 ( .A(n11), .Z(n1419) );
  BUF_X1 U26 ( .A(n7), .Z(n1440) );
  BUF_X1 U27 ( .A(n7), .Z(n1441) );
  BUF_X1 U28 ( .A(n9), .Z(n1430) );
  BUF_X1 U29 ( .A(n7), .Z(n1442) );
  BUF_X1 U30 ( .A(n7), .Z(n1439) );
  BUF_X1 U31 ( .A(n9), .Z(n1431) );
  BUF_X1 U32 ( .A(n9), .Z(n1428) );
  BUF_X1 U33 ( .A(n9), .Z(n1429) );
  BUF_X1 U34 ( .A(n9), .Z(n1427) );
  BUF_X1 U35 ( .A(n7), .Z(n1443) );
  BUF_X1 U36 ( .A(n14), .Z(n1400) );
  BUF_X1 U37 ( .A(n14), .Z(n1398) );
  BUF_X1 U38 ( .A(n14), .Z(n1399) );
  BUF_X1 U39 ( .A(n14), .Z(n1397) );
  BUF_X1 U40 ( .A(n14), .Z(n1401) );
  NOR3_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1446), .ZN(n13) );
  NOR3_X1 U42 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1445), .ZN(n12) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1446), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1446), .A2(n1445), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1445) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1446) );
  NOR3_X1 U47 ( .A1(n1446), .A2(SEL[2]), .A3(n1445), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1445), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U52 ( .A1(B[18]), .A2(n1403), .B1(A[18]), .B2(n1397), .ZN(n227) );
  AOI22_X1 U53 ( .A1(D[18]), .A2(n1415), .B1(C[18]), .B2(n1409), .ZN(n228) );
  AOI22_X1 U54 ( .A1(H[18]), .A2(n1439), .B1(G[18]), .B2(n1433), .ZN(n230) );
  NAND4_X1 U55 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U56 ( .A1(B[31]), .A2(n1405), .B1(A[31]), .B2(n1399), .ZN(n167) );
  AOI22_X1 U57 ( .A1(D[31]), .A2(n1417), .B1(C[31]), .B2(n1411), .ZN(n168) );
  AOI22_X1 U58 ( .A1(H[31]), .A2(n1441), .B1(G[31]), .B2(n1435), .ZN(n170) );
  AOI22_X1 U59 ( .A1(F[19]), .A2(n1427), .B1(E[19]), .B2(n1421), .ZN(n225) );
  NAND4_X1 U60 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U61 ( .A1(B[30]), .A2(n1404), .B1(A[30]), .B2(n1398), .ZN(n171) );
  AOI22_X1 U62 ( .A1(D[30]), .A2(n1416), .B1(C[30]), .B2(n1410), .ZN(n172) );
  AOI22_X1 U63 ( .A1(H[30]), .A2(n1440), .B1(G[30]), .B2(n1434), .ZN(n174) );
  NAND4_X1 U64 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U65 ( .A1(H[9]), .A2(n1444), .B1(G[9]), .B2(n1438), .ZN(n6) );
  AOI22_X1 U66 ( .A1(B[9]), .A2(n1408), .B1(A[9]), .B2(n1402), .ZN(n3) );
  AOI22_X1 U67 ( .A1(F[9]), .A2(n1432), .B1(E[9]), .B2(n1426), .ZN(n5) );
  NAND4_X1 U68 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U69 ( .A1(B[13]), .A2(n1403), .B1(A[13]), .B2(n1397), .ZN(n247) );
  AOI22_X1 U70 ( .A1(H[13]), .A2(n1439), .B1(G[13]), .B2(n1433), .ZN(n250) );
  AOI22_X1 U71 ( .A1(F[13]), .A2(n1427), .B1(E[13]), .B2(n1421), .ZN(n249) );
  AOI22_X1 U72 ( .A1(H[15]), .A2(n1439), .B1(G[15]), .B2(n1433), .ZN(n242) );
  NAND4_X1 U73 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U74 ( .A1(B[17]), .A2(n1403), .B1(A[17]), .B2(n1397), .ZN(n231) );
  AOI22_X1 U75 ( .A1(H[17]), .A2(n1439), .B1(G[17]), .B2(n1433), .ZN(n234) );
  AOI22_X1 U76 ( .A1(D[17]), .A2(n1415), .B1(C[17]), .B2(n1409), .ZN(n232) );
  AOI22_X1 U77 ( .A1(F[40]), .A2(n1429), .B1(E[40]), .B2(n1423), .ZN(n129) );
  AOI22_X1 U78 ( .A1(F[37]), .A2(n1429), .B1(E[37]), .B2(n1423), .ZN(n145) );
  AOI22_X1 U79 ( .A1(F[54]), .A2(n1431), .B1(E[54]), .B2(n1425), .ZN(n69) );
  AOI22_X1 U80 ( .A1(F[48]), .A2(n1430), .B1(E[48]), .B2(n1424), .ZN(n97) );
  AOI22_X1 U81 ( .A1(F[36]), .A2(n1429), .B1(E[36]), .B2(n1423), .ZN(n149) );
  AOI22_X1 U82 ( .A1(F[52]), .A2(n1430), .B1(E[52]), .B2(n1424), .ZN(n77) );
  AOI22_X1 U83 ( .A1(F[53]), .A2(n1431), .B1(E[53]), .B2(n1425), .ZN(n73) );
  AOI22_X1 U84 ( .A1(F[55]), .A2(n1431), .B1(E[55]), .B2(n1425), .ZN(n65) );
  AOI22_X1 U85 ( .A1(F[49]), .A2(n1430), .B1(E[49]), .B2(n1424), .ZN(n93) );
  AOI22_X1 U86 ( .A1(F[45]), .A2(n1430), .B1(E[45]), .B2(n1424), .ZN(n109) );
  AOI22_X1 U87 ( .A1(F[50]), .A2(n1430), .B1(E[50]), .B2(n1424), .ZN(n85) );
  AOI22_X1 U88 ( .A1(F[32]), .A2(n1429), .B1(E[32]), .B2(n1423), .ZN(n165) );
  AOI22_X1 U89 ( .A1(F[56]), .A2(n1431), .B1(E[56]), .B2(n1425), .ZN(n61) );
  AOI22_X1 U90 ( .A1(F[39]), .A2(n1429), .B1(E[39]), .B2(n1423), .ZN(n137) );
  AOI22_X1 U91 ( .A1(F[46]), .A2(n1430), .B1(E[46]), .B2(n1424), .ZN(n105) );
  AOI22_X1 U92 ( .A1(F[24]), .A2(n1428), .B1(E[24]), .B2(n1422), .ZN(n201) );
  AOI22_X1 U93 ( .A1(F[26]), .A2(n1428), .B1(E[26]), .B2(n1422), .ZN(n193) );
  AOI22_X1 U94 ( .A1(F[51]), .A2(n1430), .B1(E[51]), .B2(n1424), .ZN(n81) );
  AOI22_X1 U95 ( .A1(F[28]), .A2(n1428), .B1(E[28]), .B2(n1422), .ZN(n185) );
  AOI22_X1 U96 ( .A1(F[57]), .A2(n1431), .B1(E[57]), .B2(n1425), .ZN(n57) );
  AOI22_X1 U97 ( .A1(F[27]), .A2(n1428), .B1(E[27]), .B2(n1422), .ZN(n189) );
  AOI22_X1 U98 ( .A1(F[58]), .A2(n1431), .B1(E[58]), .B2(n1425), .ZN(n53) );
  AOI22_X1 U99 ( .A1(F[23]), .A2(n1428), .B1(E[23]), .B2(n1422), .ZN(n205) );
  AOI22_X1 U100 ( .A1(F[42]), .A2(n1430), .B1(E[42]), .B2(n1424), .ZN(n121) );
  AOI22_X1 U101 ( .A1(F[22]), .A2(n1428), .B1(E[22]), .B2(n1422), .ZN(n209) );
  AOI22_X1 U102 ( .A1(F[11]), .A2(n1427), .B1(E[11]), .B2(n1421), .ZN(n257) );
  AOI22_X1 U103 ( .A1(F[18]), .A2(n1427), .B1(E[18]), .B2(n1421), .ZN(n229) );
  AOI22_X1 U104 ( .A1(F[38]), .A2(n1429), .B1(E[38]), .B2(n1423), .ZN(n141) );
  AOI22_X1 U105 ( .A1(F[43]), .A2(n1430), .B1(E[43]), .B2(n1424), .ZN(n117) );
  AOI22_X1 U106 ( .A1(F[31]), .A2(n1429), .B1(E[31]), .B2(n1423), .ZN(n169) );
  AOI22_X1 U107 ( .A1(F[33]), .A2(n1429), .B1(E[33]), .B2(n1423), .ZN(n161) );
  AOI22_X1 U108 ( .A1(F[59]), .A2(n1431), .B1(E[59]), .B2(n1425), .ZN(n49) );
  AOI22_X1 U109 ( .A1(F[41]), .A2(n1429), .B1(E[41]), .B2(n1423), .ZN(n125) );
  AOI22_X1 U110 ( .A1(F[47]), .A2(n1430), .B1(E[47]), .B2(n1424), .ZN(n101) );
  AOI22_X1 U111 ( .A1(F[44]), .A2(n1430), .B1(E[44]), .B2(n1424), .ZN(n113) );
  AOI22_X1 U112 ( .A1(F[35]), .A2(n1429), .B1(E[35]), .B2(n1423), .ZN(n153) );
  AOI22_X1 U113 ( .A1(F[30]), .A2(n1428), .B1(E[30]), .B2(n1422), .ZN(n173) );
  AOI22_X1 U114 ( .A1(F[21]), .A2(n1428), .B1(E[21]), .B2(n1422), .ZN(n213) );
  AOI22_X1 U115 ( .A1(F[29]), .A2(n1428), .B1(E[29]), .B2(n1422), .ZN(n181) );
  AOI22_X1 U116 ( .A1(F[34]), .A2(n1429), .B1(E[34]), .B2(n1423), .ZN(n157) );
  AOI22_X1 U117 ( .A1(F[20]), .A2(n1428), .B1(E[20]), .B2(n1422), .ZN(n217) );
  AOI22_X1 U118 ( .A1(F[16]), .A2(n1427), .B1(E[16]), .B2(n1421), .ZN(n237) );
  AOI22_X1 U119 ( .A1(F[17]), .A2(n1427), .B1(E[17]), .B2(n1421), .ZN(n233) );
  AOI22_X1 U120 ( .A1(F[61]), .A2(n1431), .B1(E[61]), .B2(n1425), .ZN(n37) );
  AOI22_X1 U121 ( .A1(F[62]), .A2(n1431), .B1(E[62]), .B2(n1425), .ZN(n33) );
  AOI22_X1 U122 ( .A1(F[63]), .A2(n1431), .B1(E[63]), .B2(n1425), .ZN(n29) );
  AOI22_X1 U123 ( .A1(F[60]), .A2(n1431), .B1(E[60]), .B2(n1425), .ZN(n41) );
  AOI22_X1 U124 ( .A1(F[8]), .A2(n1432), .B1(E[8]), .B2(n1426), .ZN(n17) );
  NAND4_X1 U125 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U126 ( .A1(H[11]), .A2(n1439), .B1(G[11]), .B2(n1433), .ZN(n258) );
  AOI22_X1 U127 ( .A1(B[11]), .A2(n1403), .B1(A[11]), .B2(n1397), .ZN(n255) );
  AOI22_X1 U128 ( .A1(D[11]), .A2(n1415), .B1(C[11]), .B2(n1409), .ZN(n256) );
  AOI22_X1 U129 ( .A1(D[10]), .A2(n1415), .B1(C[10]), .B2(n1409), .ZN(n260) );
  AOI22_X1 U130 ( .A1(D[14]), .A2(n1415), .B1(C[14]), .B2(n1409), .ZN(n244) );
  AOI22_X1 U131 ( .A1(D[12]), .A2(n1415), .B1(C[12]), .B2(n1409), .ZN(n252) );
  AOI22_X1 U132 ( .A1(D[13]), .A2(n1415), .B1(C[13]), .B2(n1409), .ZN(n248) );
  AOI22_X1 U133 ( .A1(D[9]), .A2(n1420), .B1(C[9]), .B2(n1414), .ZN(n4) );
  NAND4_X1 U134 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U135 ( .A1(B[27]), .A2(n1404), .B1(A[27]), .B2(n1398), .ZN(n187) );
  AOI22_X1 U136 ( .A1(D[27]), .A2(n1416), .B1(C[27]), .B2(n1410), .ZN(n188) );
  AOI22_X1 U137 ( .A1(H[27]), .A2(n1440), .B1(G[27]), .B2(n1434), .ZN(n190) );
  NAND4_X1 U138 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U139 ( .A1(B[22]), .A2(n1404), .B1(A[22]), .B2(n1398), .ZN(n207) );
  AOI22_X1 U140 ( .A1(D[22]), .A2(n1416), .B1(C[22]), .B2(n1410), .ZN(n208) );
  AOI22_X1 U141 ( .A1(H[22]), .A2(n1440), .B1(G[22]), .B2(n1434), .ZN(n210) );
  NAND4_X1 U142 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U143 ( .A1(B[35]), .A2(n1405), .B1(A[35]), .B2(n1399), .ZN(n151) );
  AOI22_X1 U144 ( .A1(D[35]), .A2(n1417), .B1(C[35]), .B2(n1411), .ZN(n152) );
  AOI22_X1 U145 ( .A1(H[35]), .A2(n1441), .B1(G[35]), .B2(n1435), .ZN(n154) );
  NAND4_X1 U146 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U147 ( .A1(B[23]), .A2(n1404), .B1(A[23]), .B2(n1398), .ZN(n203) );
  AOI22_X1 U148 ( .A1(D[23]), .A2(n1416), .B1(C[23]), .B2(n1410), .ZN(n204) );
  AOI22_X1 U149 ( .A1(H[23]), .A2(n1440), .B1(G[23]), .B2(n1434), .ZN(n206) );
  NAND4_X1 U150 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U151 ( .A1(B[36]), .A2(n1405), .B1(A[36]), .B2(n1399), .ZN(n147) );
  AOI22_X1 U152 ( .A1(D[36]), .A2(n1417), .B1(C[36]), .B2(n1411), .ZN(n148) );
  AOI22_X1 U153 ( .A1(H[36]), .A2(n1441), .B1(G[36]), .B2(n1435), .ZN(n150) );
  NAND4_X1 U154 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U155 ( .A1(B[40]), .A2(n1405), .B1(A[40]), .B2(n1399), .ZN(n127) );
  AOI22_X1 U156 ( .A1(D[40]), .A2(n1417), .B1(C[40]), .B2(n1411), .ZN(n128) );
  AOI22_X1 U157 ( .A1(H[40]), .A2(n1441), .B1(G[40]), .B2(n1435), .ZN(n130) );
  NAND4_X1 U158 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U159 ( .A1(B[37]), .A2(n1405), .B1(A[37]), .B2(n1399), .ZN(n143) );
  AOI22_X1 U160 ( .A1(D[37]), .A2(n1417), .B1(C[37]), .B2(n1411), .ZN(n144) );
  AOI22_X1 U161 ( .A1(H[37]), .A2(n1441), .B1(G[37]), .B2(n1435), .ZN(n146) );
  NAND4_X1 U162 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U163 ( .A1(B[54]), .A2(n1407), .B1(A[54]), .B2(n1401), .ZN(n67) );
  AOI22_X1 U164 ( .A1(D[54]), .A2(n1419), .B1(C[54]), .B2(n1413), .ZN(n68) );
  AOI22_X1 U165 ( .A1(H[54]), .A2(n1443), .B1(G[54]), .B2(n1437), .ZN(n70) );
  NAND4_X1 U166 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U167 ( .A1(B[32]), .A2(n1405), .B1(A[32]), .B2(n1399), .ZN(n163) );
  AOI22_X1 U168 ( .A1(D[32]), .A2(n1417), .B1(C[32]), .B2(n1411), .ZN(n164) );
  AOI22_X1 U169 ( .A1(H[32]), .A2(n1441), .B1(G[32]), .B2(n1435), .ZN(n166) );
  NAND4_X1 U170 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U171 ( .A1(B[52]), .A2(n1406), .B1(A[52]), .B2(n1400), .ZN(n75) );
  AOI22_X1 U172 ( .A1(D[52]), .A2(n1418), .B1(C[52]), .B2(n1412), .ZN(n76) );
  AOI22_X1 U173 ( .A1(H[52]), .A2(n1442), .B1(G[52]), .B2(n1436), .ZN(n78) );
  NAND4_X1 U174 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U175 ( .A1(B[53]), .A2(n1407), .B1(A[53]), .B2(n1401), .ZN(n71) );
  AOI22_X1 U176 ( .A1(D[53]), .A2(n1419), .B1(C[53]), .B2(n1413), .ZN(n72) );
  AOI22_X1 U177 ( .A1(H[53]), .A2(n1443), .B1(G[53]), .B2(n1437), .ZN(n74) );
  NAND4_X1 U178 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U179 ( .A1(B[24]), .A2(n1404), .B1(A[24]), .B2(n1398), .ZN(n199) );
  AOI22_X1 U180 ( .A1(D[24]), .A2(n1416), .B1(C[24]), .B2(n1410), .ZN(n200) );
  AOI22_X1 U181 ( .A1(H[24]), .A2(n1440), .B1(G[24]), .B2(n1434), .ZN(n202) );
  NAND4_X1 U182 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U183 ( .A1(B[26]), .A2(n1404), .B1(A[26]), .B2(n1398), .ZN(n191) );
  AOI22_X1 U184 ( .A1(D[26]), .A2(n1416), .B1(C[26]), .B2(n1410), .ZN(n192) );
  AOI22_X1 U185 ( .A1(H[26]), .A2(n1440), .B1(G[26]), .B2(n1434), .ZN(n194) );
  NAND4_X1 U186 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U187 ( .A1(B[49]), .A2(n1406), .B1(A[49]), .B2(n1400), .ZN(n91) );
  AOI22_X1 U188 ( .A1(D[49]), .A2(n1418), .B1(C[49]), .B2(n1412), .ZN(n92) );
  AOI22_X1 U189 ( .A1(H[49]), .A2(n1442), .B1(G[49]), .B2(n1436), .ZN(n94) );
  NAND4_X1 U190 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U191 ( .A1(B[45]), .A2(n1406), .B1(A[45]), .B2(n1400), .ZN(n107) );
  AOI22_X1 U192 ( .A1(D[45]), .A2(n1418), .B1(C[45]), .B2(n1412), .ZN(n108) );
  AOI22_X1 U193 ( .A1(H[45]), .A2(n1442), .B1(G[45]), .B2(n1436), .ZN(n110) );
  NAND4_X1 U194 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U195 ( .A1(B[50]), .A2(n1406), .B1(A[50]), .B2(n1400), .ZN(n83) );
  AOI22_X1 U196 ( .A1(D[50]), .A2(n1418), .B1(C[50]), .B2(n1412), .ZN(n84) );
  AOI22_X1 U197 ( .A1(H[50]), .A2(n1442), .B1(G[50]), .B2(n1436), .ZN(n86) );
  NAND4_X1 U198 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U199 ( .A1(B[28]), .A2(n1404), .B1(A[28]), .B2(n1398), .ZN(n183) );
  AOI22_X1 U200 ( .A1(D[28]), .A2(n1416), .B1(C[28]), .B2(n1410), .ZN(n184) );
  AOI22_X1 U201 ( .A1(H[28]), .A2(n1440), .B1(G[28]), .B2(n1434), .ZN(n186) );
  NAND4_X1 U202 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U203 ( .A1(B[56]), .A2(n1407), .B1(A[56]), .B2(n1401), .ZN(n59) );
  AOI22_X1 U204 ( .A1(D[56]), .A2(n1419), .B1(C[56]), .B2(n1413), .ZN(n60) );
  AOI22_X1 U205 ( .A1(H[56]), .A2(n1443), .B1(G[56]), .B2(n1437), .ZN(n62) );
  NAND4_X1 U206 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U207 ( .A1(B[46]), .A2(n1406), .B1(A[46]), .B2(n1400), .ZN(n103) );
  AOI22_X1 U208 ( .A1(D[46]), .A2(n1418), .B1(C[46]), .B2(n1412), .ZN(n104) );
  AOI22_X1 U209 ( .A1(H[46]), .A2(n1442), .B1(G[46]), .B2(n1436), .ZN(n106) );
  NAND4_X1 U210 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U211 ( .A1(B[51]), .A2(n1406), .B1(A[51]), .B2(n1400), .ZN(n79) );
  AOI22_X1 U212 ( .A1(D[51]), .A2(n1418), .B1(C[51]), .B2(n1412), .ZN(n80) );
  AOI22_X1 U213 ( .A1(H[51]), .A2(n1442), .B1(G[51]), .B2(n1436), .ZN(n82) );
  NAND4_X1 U214 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U215 ( .A1(B[57]), .A2(n1407), .B1(A[57]), .B2(n1401), .ZN(n55) );
  AOI22_X1 U216 ( .A1(D[57]), .A2(n1419), .B1(C[57]), .B2(n1413), .ZN(n56) );
  AOI22_X1 U217 ( .A1(H[57]), .A2(n1443), .B1(G[57]), .B2(n1437), .ZN(n58) );
  NAND4_X1 U218 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U219 ( .A1(B[58]), .A2(n1407), .B1(A[58]), .B2(n1401), .ZN(n51) );
  AOI22_X1 U220 ( .A1(D[58]), .A2(n1419), .B1(C[58]), .B2(n1413), .ZN(n52) );
  AOI22_X1 U221 ( .A1(H[58]), .A2(n1443), .B1(G[58]), .B2(n1437), .ZN(n54) );
  NAND4_X1 U222 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U223 ( .A1(B[42]), .A2(n1406), .B1(A[42]), .B2(n1400), .ZN(n119) );
  AOI22_X1 U224 ( .A1(D[42]), .A2(n1418), .B1(C[42]), .B2(n1412), .ZN(n120) );
  AOI22_X1 U225 ( .A1(H[42]), .A2(n1442), .B1(G[42]), .B2(n1436), .ZN(n122) );
  NAND4_X1 U226 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U227 ( .A1(B[38]), .A2(n1405), .B1(A[38]), .B2(n1399), .ZN(n139) );
  AOI22_X1 U228 ( .A1(D[38]), .A2(n1417), .B1(C[38]), .B2(n1411), .ZN(n140) );
  AOI22_X1 U229 ( .A1(H[38]), .A2(n1441), .B1(G[38]), .B2(n1435), .ZN(n142) );
  NAND4_X1 U230 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U231 ( .A1(B[34]), .A2(n1405), .B1(A[34]), .B2(n1399), .ZN(n155) );
  AOI22_X1 U232 ( .A1(D[34]), .A2(n1417), .B1(C[34]), .B2(n1411), .ZN(n156) );
  AOI22_X1 U233 ( .A1(H[34]), .A2(n1441), .B1(G[34]), .B2(n1435), .ZN(n158) );
  NAND4_X1 U234 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U235 ( .A1(B[59]), .A2(n1407), .B1(A[59]), .B2(n1401), .ZN(n47) );
  AOI22_X1 U236 ( .A1(D[59]), .A2(n1419), .B1(C[59]), .B2(n1413), .ZN(n48) );
  AOI22_X1 U237 ( .A1(H[59]), .A2(n1443), .B1(G[59]), .B2(n1437), .ZN(n50) );
  NAND4_X1 U238 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U239 ( .A1(B[41]), .A2(n1405), .B1(A[41]), .B2(n1399), .ZN(n123) );
  AOI22_X1 U240 ( .A1(D[41]), .A2(n1417), .B1(C[41]), .B2(n1411), .ZN(n124) );
  AOI22_X1 U241 ( .A1(H[41]), .A2(n1441), .B1(G[41]), .B2(n1435), .ZN(n126) );
  NAND4_X1 U242 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U243 ( .A1(B[44]), .A2(n1406), .B1(A[44]), .B2(n1400), .ZN(n111) );
  AOI22_X1 U244 ( .A1(D[44]), .A2(n1418), .B1(C[44]), .B2(n1412), .ZN(n112) );
  AOI22_X1 U245 ( .A1(H[44]), .A2(n1442), .B1(G[44]), .B2(n1436), .ZN(n114) );
  NAND4_X1 U246 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U247 ( .A1(H[12]), .A2(n1439), .B1(G[12]), .B2(n1433), .ZN(n254) );
  AOI22_X1 U248 ( .A1(B[12]), .A2(n1403), .B1(A[12]), .B2(n1397), .ZN(n251) );
  AOI22_X1 U249 ( .A1(F[12]), .A2(n1427), .B1(E[12]), .B2(n1421), .ZN(n253) );
  NAND4_X1 U250 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U251 ( .A1(B[20]), .A2(n1404), .B1(A[20]), .B2(n1398), .ZN(n215) );
  AOI22_X1 U252 ( .A1(D[20]), .A2(n1416), .B1(C[20]), .B2(n1410), .ZN(n216) );
  AOI22_X1 U253 ( .A1(H[20]), .A2(n1440), .B1(G[20]), .B2(n1434), .ZN(n218) );
  NAND4_X1 U254 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U255 ( .A1(B[61]), .A2(n1407), .B1(A[61]), .B2(n1401), .ZN(n35) );
  AOI22_X1 U256 ( .A1(D[61]), .A2(n1419), .B1(C[61]), .B2(n1413), .ZN(n36) );
  AOI22_X1 U257 ( .A1(H[61]), .A2(n1443), .B1(G[61]), .B2(n1437), .ZN(n38) );
  NAND4_X1 U258 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U259 ( .A1(B[62]), .A2(n1407), .B1(A[62]), .B2(n1401), .ZN(n31) );
  AOI22_X1 U260 ( .A1(D[62]), .A2(n1419), .B1(C[62]), .B2(n1413), .ZN(n32) );
  AOI22_X1 U261 ( .A1(H[62]), .A2(n1443), .B1(G[62]), .B2(n1437), .ZN(n34) );
  NAND4_X1 U262 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U263 ( .A1(B[63]), .A2(n1407), .B1(A[63]), .B2(n1401), .ZN(n27) );
  AOI22_X1 U264 ( .A1(D[63]), .A2(n1419), .B1(C[63]), .B2(n1413), .ZN(n28) );
  AOI22_X1 U265 ( .A1(H[63]), .A2(n1443), .B1(G[63]), .B2(n1437), .ZN(n30) );
  NAND4_X1 U266 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U267 ( .A1(B[60]), .A2(n1407), .B1(A[60]), .B2(n1401), .ZN(n39) );
  AOI22_X1 U268 ( .A1(D[60]), .A2(n1419), .B1(C[60]), .B2(n1413), .ZN(n40) );
  AOI22_X1 U269 ( .A1(H[60]), .A2(n1443), .B1(G[60]), .B2(n1437), .ZN(n42) );
  NAND4_X1 U270 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U271 ( .A1(B[15]), .A2(n1403), .B1(A[15]), .B2(n1397), .ZN(n239) );
  AOI22_X1 U272 ( .A1(D[15]), .A2(n1415), .B1(C[15]), .B2(n1409), .ZN(n240) );
  AOI22_X1 U273 ( .A1(F[15]), .A2(n1427), .B1(E[15]), .B2(n1421), .ZN(n241) );
  NAND4_X1 U274 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U275 ( .A1(B[29]), .A2(n1404), .B1(A[29]), .B2(n1398), .ZN(n179) );
  AOI22_X1 U276 ( .A1(D[29]), .A2(n1416), .B1(C[29]), .B2(n1410), .ZN(n180) );
  AOI22_X1 U277 ( .A1(H[29]), .A2(n1440), .B1(G[29]), .B2(n1434), .ZN(n182) );
  NAND4_X1 U278 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U279 ( .A1(B[21]), .A2(n1404), .B1(A[21]), .B2(n1398), .ZN(n211) );
  AOI22_X1 U280 ( .A1(D[21]), .A2(n1416), .B1(C[21]), .B2(n1410), .ZN(n212) );
  AOI22_X1 U281 ( .A1(H[21]), .A2(n1440), .B1(G[21]), .B2(n1434), .ZN(n214) );
  NAND4_X1 U282 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U283 ( .A1(B[19]), .A2(n1403), .B1(A[19]), .B2(n1397), .ZN(n223) );
  AOI22_X1 U284 ( .A1(D[19]), .A2(n1415), .B1(C[19]), .B2(n1409), .ZN(n224) );
  AOI22_X1 U285 ( .A1(H[19]), .A2(n1439), .B1(G[19]), .B2(n1433), .ZN(n226) );
  AOI22_X1 U286 ( .A1(F[25]), .A2(n1428), .B1(E[25]), .B2(n1422), .ZN(n197) );
  NAND4_X1 U287 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U288 ( .A1(B[25]), .A2(n1404), .B1(A[25]), .B2(n1398), .ZN(n195) );
  AOI22_X1 U289 ( .A1(D[25]), .A2(n1416), .B1(C[25]), .B2(n1410), .ZN(n196) );
  AOI22_X1 U290 ( .A1(H[25]), .A2(n1440), .B1(G[25]), .B2(n1434), .ZN(n198) );
  NAND4_X1 U291 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U292 ( .A1(B[14]), .A2(n1403), .B1(A[14]), .B2(n1397), .ZN(n243) );
  AOI22_X1 U293 ( .A1(H[14]), .A2(n1439), .B1(G[14]), .B2(n1433), .ZN(n246) );
  AOI22_X1 U294 ( .A1(F[14]), .A2(n1427), .B1(E[14]), .B2(n1421), .ZN(n245) );
  NAND4_X1 U295 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U296 ( .A1(B[10]), .A2(n1403), .B1(A[10]), .B2(n1397), .ZN(n259) );
  AOI22_X1 U297 ( .A1(H[10]), .A2(n1439), .B1(G[10]), .B2(n1433), .ZN(n262) );
  AOI22_X1 U298 ( .A1(F[10]), .A2(n1427), .B1(E[10]), .B2(n1421), .ZN(n261) );
  NAND4_X1 U299 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U300 ( .A1(B[33]), .A2(n1405), .B1(A[33]), .B2(n1399), .ZN(n159) );
  AOI22_X1 U301 ( .A1(D[33]), .A2(n1417), .B1(C[33]), .B2(n1411), .ZN(n160) );
  AOI22_X1 U302 ( .A1(H[33]), .A2(n1441), .B1(G[33]), .B2(n1435), .ZN(n162) );
  NAND4_X1 U303 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U304 ( .A1(B[48]), .A2(n1406), .B1(A[48]), .B2(n1400), .ZN(n95) );
  AOI22_X1 U305 ( .A1(D[48]), .A2(n1418), .B1(C[48]), .B2(n1412), .ZN(n96) );
  AOI22_X1 U306 ( .A1(H[48]), .A2(n1442), .B1(G[48]), .B2(n1436), .ZN(n98) );
  NAND4_X1 U307 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U308 ( .A1(B[55]), .A2(n1407), .B1(A[55]), .B2(n1401), .ZN(n63) );
  AOI22_X1 U309 ( .A1(D[55]), .A2(n1419), .B1(C[55]), .B2(n1413), .ZN(n64) );
  AOI22_X1 U310 ( .A1(H[55]), .A2(n1443), .B1(G[55]), .B2(n1437), .ZN(n66) );
  NAND4_X1 U311 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U312 ( .A1(B[43]), .A2(n1406), .B1(A[43]), .B2(n1400), .ZN(n115) );
  AOI22_X1 U313 ( .A1(D[43]), .A2(n1418), .B1(C[43]), .B2(n1412), .ZN(n116) );
  AOI22_X1 U314 ( .A1(H[43]), .A2(n1442), .B1(G[43]), .B2(n1436), .ZN(n118) );
  NAND4_X1 U315 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U316 ( .A1(B[16]), .A2(n1403), .B1(A[16]), .B2(n1397), .ZN(n235) );
  AOI22_X1 U317 ( .A1(H[16]), .A2(n1439), .B1(G[16]), .B2(n1433), .ZN(n238) );
  AOI22_X1 U318 ( .A1(D[16]), .A2(n1415), .B1(C[16]), .B2(n1409), .ZN(n236) );
  NAND4_X1 U319 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U320 ( .A1(D[8]), .A2(n1420), .B1(C[8]), .B2(n1414), .ZN(n16) );
  AOI22_X1 U321 ( .A1(H[8]), .A2(n1444), .B1(G[8]), .B2(n1438), .ZN(n18) );
  AOI22_X1 U322 ( .A1(B[8]), .A2(n1408), .B1(A[8]), .B2(n1402), .ZN(n15) );
  NAND4_X1 U323 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U324 ( .A1(B[39]), .A2(n1405), .B1(A[39]), .B2(n1399), .ZN(n135) );
  AOI22_X1 U325 ( .A1(D[39]), .A2(n1417), .B1(C[39]), .B2(n1411), .ZN(n136) );
  AOI22_X1 U326 ( .A1(H[39]), .A2(n1441), .B1(G[39]), .B2(n1435), .ZN(n138) );
  NAND4_X1 U327 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U328 ( .A1(B[47]), .A2(n1406), .B1(A[47]), .B2(n1400), .ZN(n99) );
  AOI22_X1 U329 ( .A1(D[47]), .A2(n1418), .B1(C[47]), .B2(n1412), .ZN(n100) );
  AOI22_X1 U330 ( .A1(H[47]), .A2(n1442), .B1(G[47]), .B2(n1436), .ZN(n102) );
  NAND4_X1 U331 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U332 ( .A1(B[0]), .A2(n1403), .B1(A[0]), .B2(n1397), .ZN(n263) );
  AOI22_X1 U333 ( .A1(D[0]), .A2(n1415), .B1(C[0]), .B2(n1409), .ZN(n264) );
  AOI22_X1 U334 ( .A1(F[0]), .A2(n1427), .B1(E[0]), .B2(n1421), .ZN(n265) );
  NAND4_X1 U335 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U336 ( .A1(B[1]), .A2(n1403), .B1(A[1]), .B2(n1397), .ZN(n219) );
  AOI22_X1 U337 ( .A1(D[1]), .A2(n1415), .B1(C[1]), .B2(n1409), .ZN(n220) );
  AOI22_X1 U338 ( .A1(F[1]), .A2(n1427), .B1(E[1]), .B2(n1421), .ZN(n221) );
  AOI22_X1 U339 ( .A1(H[5]), .A2(n1443), .B1(G[5]), .B2(n1437), .ZN(n46) );
  AOI22_X1 U340 ( .A1(H[4]), .A2(n1442), .B1(G[4]), .B2(n1436), .ZN(n90) );
  AOI22_X1 U341 ( .A1(H[7]), .A2(n1444), .B1(G[7]), .B2(n1438), .ZN(n22) );
  AOI22_X1 U342 ( .A1(H[6]), .A2(n1444), .B1(G[6]), .B2(n1438), .ZN(n26) );
  AOI22_X1 U343 ( .A1(H[3]), .A2(n1441), .B1(G[3]), .B2(n1435), .ZN(n134) );
  AOI22_X1 U344 ( .A1(H[2]), .A2(n1440), .B1(G[2]), .B2(n1434), .ZN(n178) );
  AOI22_X1 U345 ( .A1(H[1]), .A2(n1439), .B1(G[1]), .B2(n1433), .ZN(n222) );
  NAND4_X1 U346 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U347 ( .A1(B[5]), .A2(n1407), .B1(A[5]), .B2(n1401), .ZN(n43) );
  AOI22_X1 U348 ( .A1(D[5]), .A2(n1419), .B1(C[5]), .B2(n1413), .ZN(n44) );
  AOI22_X1 U349 ( .A1(F[5]), .A2(n1431), .B1(E[5]), .B2(n1425), .ZN(n45) );
  NAND4_X1 U350 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U351 ( .A1(B[4]), .A2(n1406), .B1(A[4]), .B2(n1400), .ZN(n87) );
  AOI22_X1 U352 ( .A1(D[4]), .A2(n1418), .B1(C[4]), .B2(n1412), .ZN(n88) );
  AOI22_X1 U353 ( .A1(F[4]), .A2(n1430), .B1(E[4]), .B2(n1424), .ZN(n89) );
  NAND4_X1 U354 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U355 ( .A1(B[6]), .A2(n1408), .B1(A[6]), .B2(n1402), .ZN(n23) );
  AOI22_X1 U356 ( .A1(D[6]), .A2(n1420), .B1(C[6]), .B2(n1414), .ZN(n24) );
  AOI22_X1 U357 ( .A1(F[6]), .A2(n1432), .B1(E[6]), .B2(n1426), .ZN(n25) );
  NAND4_X1 U358 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U359 ( .A1(B[7]), .A2(n1408), .B1(A[7]), .B2(n1402), .ZN(n19) );
  AOI22_X1 U360 ( .A1(D[7]), .A2(n1420), .B1(C[7]), .B2(n1414), .ZN(n20) );
  AOI22_X1 U361 ( .A1(F[7]), .A2(n1432), .B1(E[7]), .B2(n1426), .ZN(n21) );
  NAND4_X1 U362 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U363 ( .A1(B[3]), .A2(n1405), .B1(A[3]), .B2(n1399), .ZN(n131) );
  AOI22_X1 U364 ( .A1(D[3]), .A2(n1417), .B1(C[3]), .B2(n1411), .ZN(n132) );
  AOI22_X1 U365 ( .A1(F[3]), .A2(n1429), .B1(E[3]), .B2(n1423), .ZN(n133) );
  NAND4_X1 U366 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U367 ( .A1(B[2]), .A2(n1404), .B1(A[2]), .B2(n1398), .ZN(n175) );
  AOI22_X1 U368 ( .A1(D[2]), .A2(n1416), .B1(C[2]), .B2(n1410), .ZN(n176) );
  AOI22_X1 U369 ( .A1(F[2]), .A2(n1428), .B1(E[2]), .B2(n1422), .ZN(n177) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1439), .B1(G[0]), .B2(n1433), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1402) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1408) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1414) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1420) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1426) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1432) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1438) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1444) );
endmodule


module MUX81_GENERIC_NBIT64_11 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n13), .Z(n1408) );
  BUF_X1 U2 ( .A(n13), .Z(n1407) );
  BUF_X1 U3 ( .A(n12), .Z(n1414) );
  BUF_X1 U4 ( .A(n12), .Z(n1413) );
  BUF_X1 U5 ( .A(n8), .Z(n1438) );
  BUF_X1 U6 ( .A(n8), .Z(n1437) );
  BUF_X1 U7 ( .A(n10), .Z(n1426) );
  BUF_X1 U8 ( .A(n10), .Z(n1425) );
  BUF_X1 U9 ( .A(n13), .Z(n1410) );
  BUF_X1 U10 ( .A(n13), .Z(n1409) );
  BUF_X1 U11 ( .A(n12), .Z(n1416) );
  BUF_X1 U12 ( .A(n12), .Z(n1415) );
  BUF_X1 U13 ( .A(n8), .Z(n1439) );
  BUF_X1 U14 ( .A(n8), .Z(n1440) );
  BUF_X1 U15 ( .A(n10), .Z(n1428) );
  BUF_X1 U16 ( .A(n10), .Z(n1427) );
  BUF_X1 U17 ( .A(n13), .Z(n1411) );
  BUF_X1 U18 ( .A(n12), .Z(n1417) );
  BUF_X1 U19 ( .A(n8), .Z(n1441) );
  BUF_X1 U20 ( .A(n10), .Z(n1429) );
  BUF_X1 U21 ( .A(n11), .Z(n1422) );
  BUF_X1 U22 ( .A(n11), .Z(n1420) );
  BUF_X1 U23 ( .A(n11), .Z(n1421) );
  BUF_X1 U24 ( .A(n11), .Z(n1419) );
  BUF_X1 U25 ( .A(n11), .Z(n1423) );
  BUF_X1 U26 ( .A(n7), .Z(n1444) );
  BUF_X1 U27 ( .A(n7), .Z(n1445) );
  BUF_X1 U28 ( .A(n7), .Z(n1446) );
  BUF_X1 U29 ( .A(n9), .Z(n1434) );
  BUF_X1 U30 ( .A(n7), .Z(n1443) );
  BUF_X1 U31 ( .A(n7), .Z(n1447) );
  BUF_X1 U32 ( .A(n9), .Z(n1432) );
  BUF_X1 U33 ( .A(n9), .Z(n1433) );
  BUF_X1 U34 ( .A(n9), .Z(n1431) );
  BUF_X1 U35 ( .A(n9), .Z(n1435) );
  BUF_X1 U36 ( .A(n14), .Z(n1404) );
  BUF_X1 U37 ( .A(n14), .Z(n1402) );
  BUF_X1 U38 ( .A(n14), .Z(n1403) );
  BUF_X1 U39 ( .A(n14), .Z(n1401) );
  BUF_X1 U40 ( .A(n14), .Z(n1405) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1449) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U52 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U53 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  AOI22_X1 U54 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  AOI22_X1 U55 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U56 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U57 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  NAND4_X1 U58 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U59 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U60 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  AOI22_X1 U61 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  NAND4_X1 U62 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U63 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U64 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U65 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  NAND4_X1 U66 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U67 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U68 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  AOI22_X1 U69 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  NAND4_X1 U70 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U71 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U72 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U73 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  AOI22_X1 U74 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U75 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U76 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  AOI22_X1 U77 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  AOI22_X1 U78 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U79 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U80 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U81 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  AOI22_X1 U82 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U83 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  AOI22_X1 U84 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  AOI22_X1 U85 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  AOI22_X1 U86 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  AOI22_X1 U87 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  AOI22_X1 U88 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  AOI22_X1 U89 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  AOI22_X1 U90 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  AOI22_X1 U91 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  AOI22_X1 U92 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  AOI22_X1 U93 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  AOI22_X1 U94 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  AOI22_X1 U95 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  AOI22_X1 U96 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  AOI22_X1 U97 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  AOI22_X1 U98 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  AOI22_X1 U99 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  AOI22_X1 U100 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  AOI22_X1 U101 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  AOI22_X1 U102 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  AOI22_X1 U103 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  AOI22_X1 U104 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  AOI22_X1 U105 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  AOI22_X1 U106 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  AOI22_X1 U107 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  AOI22_X1 U108 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  AOI22_X1 U109 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  AOI22_X1 U110 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  AOI22_X1 U111 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  AOI22_X1 U112 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  AOI22_X1 U113 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  AOI22_X1 U114 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  AOI22_X1 U115 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  AOI22_X1 U116 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  AOI22_X1 U117 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  NAND4_X1 U118 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U119 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U120 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  AOI22_X1 U121 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  NAND4_X1 U122 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U123 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  AOI22_X1 U124 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U125 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  NAND4_X1 U126 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U127 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U128 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U129 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U130 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U131 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U132 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  AOI22_X1 U133 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  AOI22_X1 U134 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  AOI22_X1 U135 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U136 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U137 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U138 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U139 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  NAND4_X1 U140 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U141 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U142 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U143 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  AOI22_X1 U144 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  AOI22_X1 U145 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U146 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U147 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  NAND4_X1 U148 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U149 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U150 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U151 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U152 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  AOI22_X1 U153 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  NAND4_X1 U154 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U155 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U156 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U157 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  NAND4_X1 U158 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U159 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U160 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  AOI22_X1 U161 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  NAND4_X1 U162 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U163 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U164 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U165 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U166 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U167 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  AOI22_X1 U168 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  AOI22_X1 U169 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  NAND4_X1 U170 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U171 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  AOI22_X1 U172 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  AOI22_X1 U173 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  NAND4_X1 U174 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U175 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U176 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  AOI22_X1 U177 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  NAND4_X1 U178 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U179 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U180 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  AOI22_X1 U181 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  NAND4_X1 U182 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U183 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U184 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  AOI22_X1 U185 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  NAND4_X1 U186 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U187 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U188 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U189 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  NAND4_X1 U190 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U191 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U192 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U193 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  NAND4_X1 U194 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U195 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U196 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U197 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  NAND4_X1 U198 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U199 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U200 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U201 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  NAND4_X1 U202 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U203 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U204 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U205 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  NAND4_X1 U206 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U207 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U208 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U209 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  NAND4_X1 U210 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U211 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U212 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U213 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  NAND4_X1 U214 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U215 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U216 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U217 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  NAND4_X1 U218 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U219 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U220 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U221 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  NAND4_X1 U222 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U223 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U224 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U225 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  NAND4_X1 U226 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U227 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U228 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U229 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  NAND4_X1 U230 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U231 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U232 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U233 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  NAND4_X1 U234 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U235 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U236 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U237 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  NAND4_X1 U238 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U239 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U240 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U241 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  NAND4_X1 U242 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U243 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U244 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U245 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  NAND4_X1 U246 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U247 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U248 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U249 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  NAND4_X1 U250 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U251 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U252 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U253 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  NAND4_X1 U254 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U255 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U256 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U257 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U258 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U259 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U260 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  AOI22_X1 U261 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  NAND4_X1 U262 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U263 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U264 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  AOI22_X1 U265 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  NAND4_X1 U266 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U267 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  AOI22_X1 U268 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  AOI22_X1 U269 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  NAND4_X1 U270 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U271 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U272 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U273 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  NAND4_X1 U274 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U275 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U276 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  AOI22_X1 U277 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  AOI22_X1 U278 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  AOI22_X1 U279 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  NAND4_X1 U280 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U281 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U282 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U283 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  NAND4_X1 U284 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U285 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U286 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U287 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  NAND4_X1 U288 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U289 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U290 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U291 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  NAND4_X1 U292 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U293 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U294 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U295 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  NAND4_X1 U296 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U297 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U298 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U299 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  NAND4_X1 U300 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U301 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U302 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U303 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  NAND4_X1 U304 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U305 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U306 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U307 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  NAND4_X1 U308 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U309 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U310 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U311 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  NAND4_X1 U312 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U313 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U314 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U315 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  NAND4_X1 U316 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U317 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U318 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U319 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  NAND4_X1 U320 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U321 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U322 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U323 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U324 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U325 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U326 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U327 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U328 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U329 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U330 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U331 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U332 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U333 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U334 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U335 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U336 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U337 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U338 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U339 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U340 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U341 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U342 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U343 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U344 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U345 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U346 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U347 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U348 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U349 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U350 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U351 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U352 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U353 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U354 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U355 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U356 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U357 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U358 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U359 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U360 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U361 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U362 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U363 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U364 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U365 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U366 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U367 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U368 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U369 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  NAND4_X1 U370 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_10 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n13), .Z(n1407) );
  BUF_X1 U2 ( .A(n12), .Z(n1413) );
  BUF_X1 U3 ( .A(n8), .Z(n1437) );
  BUF_X1 U4 ( .A(n10), .Z(n1425) );
  BUF_X1 U5 ( .A(n13), .Z(n1408) );
  BUF_X1 U6 ( .A(n13), .Z(n1409) );
  BUF_X1 U7 ( .A(n12), .Z(n1416) );
  BUF_X1 U8 ( .A(n12), .Z(n1414) );
  BUF_X1 U9 ( .A(n12), .Z(n1415) );
  BUF_X1 U10 ( .A(n8), .Z(n1438) );
  BUF_X1 U11 ( .A(n8), .Z(n1439) );
  BUF_X1 U12 ( .A(n10), .Z(n1428) );
  BUF_X1 U13 ( .A(n10), .Z(n1426) );
  BUF_X1 U14 ( .A(n10), .Z(n1427) );
  BUF_X1 U15 ( .A(n13), .Z(n1410) );
  BUF_X1 U16 ( .A(n13), .Z(n1411) );
  BUF_X1 U17 ( .A(n12), .Z(n1417) );
  BUF_X1 U18 ( .A(n8), .Z(n1440) );
  BUF_X1 U19 ( .A(n8), .Z(n1441) );
  BUF_X1 U20 ( .A(n10), .Z(n1429) );
  BUF_X1 U21 ( .A(n11), .Z(n1422) );
  BUF_X1 U22 ( .A(n11), .Z(n1423) );
  BUF_X1 U23 ( .A(n11), .Z(n1420) );
  BUF_X1 U24 ( .A(n11), .Z(n1421) );
  BUF_X1 U25 ( .A(n11), .Z(n1419) );
  BUF_X1 U26 ( .A(n7), .Z(n1444) );
  BUF_X1 U27 ( .A(n7), .Z(n1445) );
  BUF_X1 U28 ( .A(n7), .Z(n1446) );
  BUF_X1 U29 ( .A(n9), .Z(n1434) );
  BUF_X1 U30 ( .A(n7), .Z(n1443) );
  BUF_X1 U31 ( .A(n7), .Z(n1447) );
  BUF_X1 U32 ( .A(n9), .Z(n1435) );
  BUF_X1 U33 ( .A(n9), .Z(n1432) );
  BUF_X1 U34 ( .A(n9), .Z(n1433) );
  BUF_X1 U35 ( .A(n9), .Z(n1431) );
  BUF_X1 U36 ( .A(n14), .Z(n1404) );
  BUF_X1 U37 ( .A(n14), .Z(n1405) );
  BUF_X1 U38 ( .A(n14), .Z(n1402) );
  BUF_X1 U39 ( .A(n14), .Z(n1403) );
  BUF_X1 U40 ( .A(n14), .Z(n1401) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1449) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U52 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U53 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  AOI22_X1 U54 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  AOI22_X1 U55 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  AOI22_X1 U56 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U57 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  NAND4_X1 U58 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U59 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  AOI22_X1 U60 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U61 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  NAND4_X1 U62 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U63 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  AOI22_X1 U64 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  AOI22_X1 U65 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  NAND4_X1 U66 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U67 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U68 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U69 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  NAND4_X1 U70 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U71 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U72 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  AOI22_X1 U73 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  NAND4_X1 U74 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U75 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U76 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U77 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U78 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U79 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U80 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U81 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  NAND4_X1 U82 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U83 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U84 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U85 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  NAND4_X1 U86 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U87 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U88 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  AOI22_X1 U89 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  AOI22_X1 U90 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U91 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U92 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  AOI22_X1 U93 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U94 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  AOI22_X1 U95 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  AOI22_X1 U96 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  AOI22_X1 U97 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  AOI22_X1 U98 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  AOI22_X1 U99 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  AOI22_X1 U100 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  AOI22_X1 U101 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  AOI22_X1 U102 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  AOI22_X1 U103 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  AOI22_X1 U104 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  AOI22_X1 U105 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  AOI22_X1 U106 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  AOI22_X1 U107 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  AOI22_X1 U108 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  AOI22_X1 U109 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  AOI22_X1 U110 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  AOI22_X1 U111 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  AOI22_X1 U112 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  AOI22_X1 U113 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  AOI22_X1 U114 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  AOI22_X1 U115 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  AOI22_X1 U116 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  AOI22_X1 U117 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  AOI22_X1 U118 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  AOI22_X1 U119 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  AOI22_X1 U120 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  AOI22_X1 U121 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  AOI22_X1 U122 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  AOI22_X1 U123 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  AOI22_X1 U124 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  AOI22_X1 U125 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  AOI22_X1 U126 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  AOI22_X1 U127 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  AOI22_X1 U128 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  AOI22_X1 U129 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  AOI22_X1 U130 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  AOI22_X1 U131 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  AOI22_X1 U132 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  AOI22_X1 U133 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  AOI22_X1 U134 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  AOI22_X1 U135 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  NAND4_X1 U136 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U137 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  AOI22_X1 U138 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  AOI22_X1 U139 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  AOI22_X1 U140 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U141 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  NAND4_X1 U142 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U143 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U144 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  AOI22_X1 U145 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  NAND4_X1 U146 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U147 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U148 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U149 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  NAND4_X1 U150 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U151 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  AOI22_X1 U152 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U153 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  NAND4_X1 U154 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U155 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  AOI22_X1 U156 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  AOI22_X1 U157 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  NAND4_X1 U158 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U159 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U160 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  AOI22_X1 U161 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  NAND4_X1 U162 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U163 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U164 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  AOI22_X1 U165 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  NAND4_X1 U166 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U167 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U168 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  AOI22_X1 U169 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  NAND4_X1 U170 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U171 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U172 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U173 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  NAND4_X1 U174 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U175 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U176 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U177 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  NAND4_X1 U178 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U179 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U180 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U181 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  NAND4_X1 U182 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U183 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U184 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U185 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  NAND4_X1 U186 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U187 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U188 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U189 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  NAND4_X1 U190 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U191 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U192 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U193 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  NAND4_X1 U194 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U195 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U196 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U197 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  NAND4_X1 U198 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U199 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U200 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U201 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  NAND4_X1 U202 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U203 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U204 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U205 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  NAND4_X1 U206 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U207 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U208 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U209 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  NAND4_X1 U210 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U211 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U212 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U213 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  NAND4_X1 U214 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U215 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U216 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U217 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  NAND4_X1 U218 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U219 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U220 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U221 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  NAND4_X1 U222 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U223 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U224 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U225 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  NAND4_X1 U226 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U227 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U228 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U229 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  NAND4_X1 U230 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U231 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U232 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U233 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  NAND4_X1 U234 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U235 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U236 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U237 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  NAND4_X1 U238 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U239 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U240 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U241 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  NAND4_X1 U242 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U243 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U244 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U245 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  NAND4_X1 U246 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U247 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U248 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U249 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  NAND4_X1 U250 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U251 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U252 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U253 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  NAND4_X1 U254 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U255 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U256 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U257 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  NAND4_X1 U258 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U259 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U260 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U261 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  NAND4_X1 U262 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U263 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U264 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  AOI22_X1 U265 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  NAND4_X1 U266 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U267 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U268 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U269 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  NAND4_X1 U270 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U271 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U272 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U273 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  NAND4_X1 U274 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U275 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U276 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U277 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  NAND4_X1 U278 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U279 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U280 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U281 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  NAND4_X1 U282 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U283 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U284 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U285 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  NAND4_X1 U286 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U287 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U288 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U289 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  NAND4_X1 U290 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U291 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U292 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U293 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U294 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U295 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U296 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  AOI22_X1 U297 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  NAND4_X1 U298 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U299 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U300 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U301 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  NAND4_X1 U302 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U303 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U304 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U305 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  NAND4_X1 U306 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U307 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U308 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U309 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  AOI22_X1 U310 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  NAND4_X1 U311 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U312 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U313 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U314 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U315 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U316 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U317 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U318 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U319 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U320 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U321 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U322 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U323 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U324 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U325 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U326 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U327 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U328 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U329 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U330 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U331 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U332 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U333 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U334 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U335 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U336 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U337 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U338 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U339 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U340 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U341 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U342 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U343 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U344 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U345 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U346 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U347 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U348 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U349 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U350 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U351 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U352 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U353 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U354 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U355 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U356 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U357 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U358 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U359 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U360 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U361 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U362 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U363 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U364 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U365 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_9 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n12), .Z(n1413) );
  BUF_X1 U2 ( .A(n10), .Z(n1425) );
  BUF_X1 U3 ( .A(n13), .Z(n1408) );
  BUF_X1 U4 ( .A(n13), .Z(n1409) );
  BUF_X1 U5 ( .A(n13), .Z(n1407) );
  BUF_X1 U6 ( .A(n12), .Z(n1414) );
  BUF_X1 U7 ( .A(n12), .Z(n1415) );
  BUF_X1 U8 ( .A(n8), .Z(n1438) );
  BUF_X1 U9 ( .A(n8), .Z(n1439) );
  BUF_X1 U10 ( .A(n8), .Z(n1437) );
  BUF_X1 U11 ( .A(n10), .Z(n1426) );
  BUF_X1 U12 ( .A(n10), .Z(n1427) );
  BUF_X1 U13 ( .A(n13), .Z(n1410) );
  BUF_X1 U14 ( .A(n13), .Z(n1411) );
  BUF_X1 U15 ( .A(n12), .Z(n1416) );
  BUF_X1 U16 ( .A(n12), .Z(n1417) );
  BUF_X1 U17 ( .A(n10), .Z(n1428) );
  BUF_X1 U18 ( .A(n8), .Z(n1440) );
  BUF_X1 U19 ( .A(n10), .Z(n1429) );
  BUF_X1 U20 ( .A(n8), .Z(n1441) );
  BUF_X1 U21 ( .A(n11), .Z(n1422) );
  BUF_X1 U22 ( .A(n11), .Z(n1423) );
  BUF_X1 U23 ( .A(n11), .Z(n1420) );
  BUF_X1 U24 ( .A(n11), .Z(n1421) );
  BUF_X1 U25 ( .A(n11), .Z(n1419) );
  BUF_X1 U26 ( .A(n7), .Z(n1444) );
  BUF_X1 U27 ( .A(n7), .Z(n1445) );
  BUF_X1 U28 ( .A(n9), .Z(n1434) );
  BUF_X1 U29 ( .A(n7), .Z(n1446) );
  BUF_X1 U30 ( .A(n7), .Z(n1443) );
  BUF_X1 U31 ( .A(n9), .Z(n1435) );
  BUF_X1 U32 ( .A(n7), .Z(n1447) );
  BUF_X1 U33 ( .A(n9), .Z(n1432) );
  BUF_X1 U34 ( .A(n9), .Z(n1433) );
  BUF_X1 U35 ( .A(n9), .Z(n1431) );
  BUF_X1 U36 ( .A(n14), .Z(n1404) );
  BUF_X1 U37 ( .A(n14), .Z(n1405) );
  BUF_X1 U38 ( .A(n14), .Z(n1402) );
  BUF_X1 U39 ( .A(n14), .Z(n1403) );
  BUF_X1 U40 ( .A(n14), .Z(n1401) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  AND3_X1 U42 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U43 ( .A(SEL[1]), .ZN(n1449) );
  NOR3_X1 U44 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U45 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  AOI22_X1 U51 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  AOI22_X1 U52 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  NAND4_X1 U53 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U54 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  AOI22_X1 U55 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U56 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  NAND4_X1 U57 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U58 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  AOI22_X1 U59 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U60 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  NAND4_X1 U61 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U62 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U63 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  AOI22_X1 U64 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  NAND4_X1 U65 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U66 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U67 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  AOI22_X1 U68 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  NAND4_X1 U69 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U70 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U71 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U72 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  NAND4_X1 U73 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U74 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U75 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U76 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  AOI22_X1 U77 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  AOI22_X1 U78 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  AOI22_X1 U79 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  AOI22_X1 U80 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  AOI22_X1 U81 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  AOI22_X1 U82 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  AOI22_X1 U83 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  AOI22_X1 U84 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  AOI22_X1 U85 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  AOI22_X1 U86 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  AOI22_X1 U87 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  AOI22_X1 U88 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  AOI22_X1 U89 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  AOI22_X1 U90 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  AOI22_X1 U91 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  AOI22_X1 U92 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  AOI22_X1 U93 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  AOI22_X1 U94 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  AOI22_X1 U95 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  AOI22_X1 U96 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  AOI22_X1 U97 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  AOI22_X1 U98 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  AOI22_X1 U99 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  AOI22_X1 U100 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  AOI22_X1 U101 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  AOI22_X1 U102 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  AOI22_X1 U103 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  AOI22_X1 U104 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  NAND4_X1 U105 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U106 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U107 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U108 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  AOI22_X1 U109 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  AOI22_X1 U110 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  NAND4_X1 U111 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U112 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  AOI22_X1 U113 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  AOI22_X1 U114 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  NAND4_X1 U115 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U116 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U117 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U118 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  NAND4_X1 U119 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U120 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U121 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  AOI22_X1 U122 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  NAND4_X1 U123 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U124 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U125 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U126 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  NAND4_X1 U127 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U128 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U129 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U130 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  NAND4_X1 U131 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U132 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U133 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U134 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  NAND4_X1 U135 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U136 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U137 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U138 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  NAND4_X1 U139 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U140 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U141 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U142 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  NAND4_X1 U143 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U144 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U145 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U146 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  NAND4_X1 U147 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U148 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U149 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  AOI22_X1 U150 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  NAND4_X1 U151 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U152 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U153 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U154 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  NAND4_X1 U155 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U156 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U157 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U158 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  NAND4_X1 U159 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U160 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U161 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U162 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  NAND4_X1 U163 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U164 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U165 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U166 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  NAND4_X1 U167 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U168 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U169 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U170 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  NAND4_X1 U171 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U172 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U173 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U174 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  NAND4_X1 U175 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U176 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U177 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U178 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  NAND4_X1 U179 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U180 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U181 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U182 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  NAND4_X1 U183 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U184 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  AOI22_X1 U185 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U186 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  NAND4_X1 U187 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U188 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  AOI22_X1 U189 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U190 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  NAND4_X1 U191 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U192 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U193 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U194 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  NAND4_X1 U195 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U196 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U197 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U198 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  NAND4_X1 U199 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U200 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U201 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  AOI22_X1 U202 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  NAND4_X1 U203 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U204 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U205 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U206 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  NAND4_X1 U207 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U208 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U209 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U210 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  NAND4_X1 U211 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U212 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U213 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  AOI22_X1 U214 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  NAND4_X1 U215 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U216 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U217 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U218 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  AOI22_X1 U219 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  AOI22_X1 U220 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  AOI22_X1 U221 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  AOI22_X1 U222 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  AOI22_X1 U223 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  AOI22_X1 U224 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  AOI22_X1 U225 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  AOI22_X1 U226 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  AOI22_X1 U227 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  AOI22_X1 U228 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  AOI22_X1 U229 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  AOI22_X1 U230 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  AOI22_X1 U231 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  AOI22_X1 U232 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  AOI22_X1 U233 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  AOI22_X1 U234 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  AOI22_X1 U235 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  NAND4_X1 U236 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U237 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U238 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U239 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  NAND4_X1 U240 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U241 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U242 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U243 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  NAND4_X1 U244 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U245 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U246 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U247 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  NAND4_X1 U248 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U249 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U250 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U251 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  NAND4_X1 U252 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U253 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U254 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U255 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  NAND4_X1 U256 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U257 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U258 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U259 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  NAND4_X1 U260 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U261 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U262 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U263 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  NAND4_X1 U264 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U265 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U266 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U267 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  NAND4_X1 U268 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U269 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U270 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U271 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  NAND4_X1 U272 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U273 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U274 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U275 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  NAND4_X1 U276 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U277 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U278 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U279 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  NAND4_X1 U280 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U281 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U282 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U283 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  NAND4_X1 U284 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U285 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U286 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U287 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  NAND4_X1 U288 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U289 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U290 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U291 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  NAND4_X1 U292 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U293 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U294 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U295 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  NAND4_X1 U296 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U297 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U298 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U299 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  AOI22_X1 U300 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U301 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U302 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U303 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U304 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U305 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U306 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U307 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U308 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U309 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U310 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U311 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U312 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U313 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U314 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U315 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U316 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U317 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U318 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U319 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U320 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U321 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U322 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U323 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U324 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U325 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U326 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U327 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U328 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U329 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U330 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U331 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U332 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U333 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U334 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U335 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U336 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U337 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U338 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U339 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U340 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U341 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U342 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U343 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  AOI22_X1 U344 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  AOI22_X1 U345 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  NAND4_X1 U346 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U347 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U348 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U349 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U350 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U351 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U352 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U353 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U354 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U355 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U356 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U357 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U358 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U359 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U360 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U361 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U362 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U363 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U364 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U365 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_8 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446;

  BUF_X1 U1 ( .A(n13), .Z(n1404) );
  BUF_X1 U2 ( .A(n13), .Z(n1403) );
  BUF_X1 U3 ( .A(n12), .Z(n1410) );
  BUF_X1 U4 ( .A(n12), .Z(n1411) );
  BUF_X1 U5 ( .A(n12), .Z(n1409) );
  BUF_X1 U6 ( .A(n8), .Z(n1433) );
  BUF_X1 U7 ( .A(n8), .Z(n1434) );
  BUF_X1 U8 ( .A(n10), .Z(n1422) );
  BUF_X1 U9 ( .A(n10), .Z(n1423) );
  BUF_X1 U10 ( .A(n10), .Z(n1421) );
  BUF_X1 U11 ( .A(n13), .Z(n1406) );
  BUF_X1 U12 ( .A(n13), .Z(n1405) );
  BUF_X1 U13 ( .A(n12), .Z(n1412) );
  BUF_X1 U14 ( .A(n8), .Z(n1435) );
  BUF_X1 U15 ( .A(n10), .Z(n1424) );
  BUF_X1 U16 ( .A(n8), .Z(n1436) );
  BUF_X1 U17 ( .A(n13), .Z(n1407) );
  BUF_X1 U18 ( .A(n12), .Z(n1413) );
  BUF_X1 U19 ( .A(n10), .Z(n1425) );
  BUF_X1 U20 ( .A(n8), .Z(n1437) );
  BUF_X1 U21 ( .A(n11), .Z(n1418) );
  BUF_X1 U22 ( .A(n11), .Z(n1419) );
  BUF_X1 U23 ( .A(n11), .Z(n1416) );
  BUF_X1 U24 ( .A(n11), .Z(n1417) );
  BUF_X1 U25 ( .A(n11), .Z(n1415) );
  BUF_X1 U26 ( .A(n7), .Z(n1439) );
  BUF_X1 U27 ( .A(n7), .Z(n1440) );
  BUF_X1 U28 ( .A(n7), .Z(n1441) );
  BUF_X1 U29 ( .A(n9), .Z(n1430) );
  BUF_X1 U30 ( .A(n7), .Z(n1442) );
  BUF_X1 U31 ( .A(n9), .Z(n1431) );
  BUF_X1 U32 ( .A(n7), .Z(n1443) );
  BUF_X1 U33 ( .A(n9), .Z(n1428) );
  BUF_X1 U34 ( .A(n9), .Z(n1429) );
  BUF_X1 U35 ( .A(n9), .Z(n1427) );
  BUF_X1 U36 ( .A(n14), .Z(n1400) );
  BUF_X1 U37 ( .A(n14), .Z(n1401) );
  BUF_X1 U38 ( .A(n14), .Z(n1398) );
  BUF_X1 U39 ( .A(n14), .Z(n1399) );
  BUF_X1 U40 ( .A(n14), .Z(n1397) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1445), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1446), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1446), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1446), .A2(n1445), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1445) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1446) );
  NOR3_X1 U47 ( .A1(n1446), .A2(SEL[2]), .A3(n1445), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1445), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U52 ( .A1(B[24]), .A2(n1404), .B1(A[24]), .B2(n1398), .ZN(n199) );
  AOI22_X1 U53 ( .A1(D[24]), .A2(n1416), .B1(C[24]), .B2(n1410), .ZN(n200) );
  AOI22_X1 U54 ( .A1(H[24]), .A2(n1440), .B1(G[24]), .B2(n1434), .ZN(n202) );
  NAND4_X1 U55 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U56 ( .A1(B[26]), .A2(n1404), .B1(A[26]), .B2(n1398), .ZN(n191) );
  AOI22_X1 U57 ( .A1(D[26]), .A2(n1416), .B1(C[26]), .B2(n1410), .ZN(n192) );
  AOI22_X1 U58 ( .A1(H[26]), .A2(n1440), .B1(G[26]), .B2(n1434), .ZN(n194) );
  AOI22_X1 U59 ( .A1(F[62]), .A2(n1431), .B1(E[62]), .B2(n1425), .ZN(n33) );
  AOI22_X1 U60 ( .A1(F[61]), .A2(n1431), .B1(E[61]), .B2(n1425), .ZN(n37) );
  NAND4_X1 U61 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U62 ( .A1(B[37]), .A2(n1405), .B1(A[37]), .B2(n1399), .ZN(n143) );
  AOI22_X1 U63 ( .A1(D[37]), .A2(n1417), .B1(C[37]), .B2(n1411), .ZN(n144) );
  AOI22_X1 U64 ( .A1(H[37]), .A2(n1441), .B1(G[37]), .B2(n1435), .ZN(n146) );
  NAND4_X1 U65 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U66 ( .A1(H[19]), .A2(n1439), .B1(G[19]), .B2(n1433), .ZN(n226) );
  AOI22_X1 U67 ( .A1(B[19]), .A2(n1403), .B1(A[19]), .B2(n1397), .ZN(n223) );
  AOI22_X1 U68 ( .A1(F[19]), .A2(n1427), .B1(E[19]), .B2(n1421), .ZN(n225) );
  NAND4_X1 U69 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U70 ( .A1(B[46]), .A2(n1406), .B1(A[46]), .B2(n1400), .ZN(n103) );
  AOI22_X1 U71 ( .A1(D[46]), .A2(n1418), .B1(C[46]), .B2(n1412), .ZN(n104) );
  AOI22_X1 U72 ( .A1(H[46]), .A2(n1442), .B1(G[46]), .B2(n1436), .ZN(n106) );
  NAND4_X1 U73 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U74 ( .A1(B[40]), .A2(n1405), .B1(A[40]), .B2(n1399), .ZN(n127) );
  AOI22_X1 U75 ( .A1(D[40]), .A2(n1417), .B1(C[40]), .B2(n1411), .ZN(n128) );
  AOI22_X1 U76 ( .A1(H[40]), .A2(n1441), .B1(G[40]), .B2(n1435), .ZN(n130) );
  NAND4_X1 U77 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U78 ( .A1(B[23]), .A2(n1404), .B1(A[23]), .B2(n1398), .ZN(n203) );
  AOI22_X1 U79 ( .A1(D[23]), .A2(n1416), .B1(C[23]), .B2(n1410), .ZN(n204) );
  AOI22_X1 U80 ( .A1(H[23]), .A2(n1440), .B1(G[23]), .B2(n1434), .ZN(n206) );
  NAND4_X1 U81 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U82 ( .A1(B[35]), .A2(n1405), .B1(A[35]), .B2(n1399), .ZN(n151) );
  AOI22_X1 U83 ( .A1(D[35]), .A2(n1417), .B1(C[35]), .B2(n1411), .ZN(n152) );
  AOI22_X1 U84 ( .A1(H[35]), .A2(n1441), .B1(G[35]), .B2(n1435), .ZN(n154) );
  NAND4_X1 U85 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U86 ( .A1(B[47]), .A2(n1406), .B1(A[47]), .B2(n1400), .ZN(n99) );
  AOI22_X1 U87 ( .A1(D[47]), .A2(n1418), .B1(C[47]), .B2(n1412), .ZN(n100) );
  AOI22_X1 U88 ( .A1(H[47]), .A2(n1442), .B1(G[47]), .B2(n1436), .ZN(n102) );
  NAND4_X1 U89 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U90 ( .A1(B[34]), .A2(n1405), .B1(A[34]), .B2(n1399), .ZN(n155) );
  AOI22_X1 U91 ( .A1(D[34]), .A2(n1417), .B1(C[34]), .B2(n1411), .ZN(n156) );
  AOI22_X1 U92 ( .A1(H[34]), .A2(n1441), .B1(G[34]), .B2(n1435), .ZN(n158) );
  NAND4_X1 U93 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U94 ( .A1(B[27]), .A2(n1404), .B1(A[27]), .B2(n1398), .ZN(n187) );
  AOI22_X1 U95 ( .A1(D[27]), .A2(n1416), .B1(C[27]), .B2(n1410), .ZN(n188) );
  AOI22_X1 U96 ( .A1(H[27]), .A2(n1440), .B1(G[27]), .B2(n1434), .ZN(n190) );
  AOI22_X1 U97 ( .A1(F[16]), .A2(n1427), .B1(E[16]), .B2(n1421), .ZN(n237) );
  AOI22_X1 U98 ( .A1(F[23]), .A2(n1428), .B1(E[23]), .B2(n1422), .ZN(n205) );
  AOI22_X1 U99 ( .A1(F[25]), .A2(n1428), .B1(E[25]), .B2(n1422), .ZN(n197) );
  AOI22_X1 U100 ( .A1(F[21]), .A2(n1428), .B1(E[21]), .B2(n1422), .ZN(n213) );
  AOI22_X1 U101 ( .A1(F[20]), .A2(n1428), .B1(E[20]), .B2(n1422), .ZN(n217) );
  AOI22_X1 U102 ( .A1(F[22]), .A2(n1428), .B1(E[22]), .B2(n1422), .ZN(n209) );
  AOI22_X1 U103 ( .A1(F[27]), .A2(n1428), .B1(E[27]), .B2(n1422), .ZN(n189) );
  AOI22_X1 U104 ( .A1(F[26]), .A2(n1428), .B1(E[26]), .B2(n1422), .ZN(n193) );
  AOI22_X1 U105 ( .A1(F[24]), .A2(n1428), .B1(E[24]), .B2(n1422), .ZN(n201) );
  AOI22_X1 U106 ( .A1(F[31]), .A2(n1429), .B1(E[31]), .B2(n1423), .ZN(n169) );
  AOI22_X1 U107 ( .A1(F[28]), .A2(n1428), .B1(E[28]), .B2(n1422), .ZN(n185) );
  AOI22_X1 U108 ( .A1(F[29]), .A2(n1428), .B1(E[29]), .B2(n1422), .ZN(n181) );
  AOI22_X1 U109 ( .A1(F[30]), .A2(n1428), .B1(E[30]), .B2(n1422), .ZN(n173) );
  AOI22_X1 U110 ( .A1(F[33]), .A2(n1429), .B1(E[33]), .B2(n1423), .ZN(n161) );
  AOI22_X1 U111 ( .A1(F[35]), .A2(n1429), .B1(E[35]), .B2(n1423), .ZN(n153) );
  AOI22_X1 U112 ( .A1(F[34]), .A2(n1429), .B1(E[34]), .B2(n1423), .ZN(n157) );
  AOI22_X1 U113 ( .A1(F[32]), .A2(n1429), .B1(E[32]), .B2(n1423), .ZN(n165) );
  AOI22_X1 U114 ( .A1(F[38]), .A2(n1429), .B1(E[38]), .B2(n1423), .ZN(n141) );
  AOI22_X1 U115 ( .A1(F[39]), .A2(n1429), .B1(E[39]), .B2(n1423), .ZN(n137) );
  AOI22_X1 U116 ( .A1(F[36]), .A2(n1429), .B1(E[36]), .B2(n1423), .ZN(n149) );
  AOI22_X1 U117 ( .A1(F[41]), .A2(n1429), .B1(E[41]), .B2(n1423), .ZN(n125) );
  AOI22_X1 U118 ( .A1(F[43]), .A2(n1430), .B1(E[43]), .B2(n1424), .ZN(n117) );
  AOI22_X1 U119 ( .A1(F[42]), .A2(n1430), .B1(E[42]), .B2(n1424), .ZN(n121) );
  AOI22_X1 U120 ( .A1(F[37]), .A2(n1429), .B1(E[37]), .B2(n1423), .ZN(n145) );
  AOI22_X1 U121 ( .A1(F[45]), .A2(n1430), .B1(E[45]), .B2(n1424), .ZN(n109) );
  AOI22_X1 U122 ( .A1(F[46]), .A2(n1430), .B1(E[46]), .B2(n1424), .ZN(n105) );
  AOI22_X1 U123 ( .A1(F[47]), .A2(n1430), .B1(E[47]), .B2(n1424), .ZN(n101) );
  AOI22_X1 U124 ( .A1(F[49]), .A2(n1430), .B1(E[49]), .B2(n1424), .ZN(n93) );
  AOI22_X1 U125 ( .A1(F[50]), .A2(n1430), .B1(E[50]), .B2(n1424), .ZN(n85) );
  AOI22_X1 U126 ( .A1(F[48]), .A2(n1430), .B1(E[48]), .B2(n1424), .ZN(n97) );
  AOI22_X1 U127 ( .A1(F[51]), .A2(n1430), .B1(E[51]), .B2(n1424), .ZN(n81) );
  AOI22_X1 U128 ( .A1(F[55]), .A2(n1431), .B1(E[55]), .B2(n1425), .ZN(n65) );
  AOI22_X1 U129 ( .A1(F[53]), .A2(n1431), .B1(E[53]), .B2(n1425), .ZN(n73) );
  AOI22_X1 U130 ( .A1(F[52]), .A2(n1430), .B1(E[52]), .B2(n1424), .ZN(n77) );
  AOI22_X1 U131 ( .A1(F[54]), .A2(n1431), .B1(E[54]), .B2(n1425), .ZN(n69) );
  AOI22_X1 U132 ( .A1(F[56]), .A2(n1431), .B1(E[56]), .B2(n1425), .ZN(n61) );
  AOI22_X1 U133 ( .A1(F[57]), .A2(n1431), .B1(E[57]), .B2(n1425), .ZN(n57) );
  AOI22_X1 U134 ( .A1(F[59]), .A2(n1431), .B1(E[59]), .B2(n1425), .ZN(n49) );
  AOI22_X1 U135 ( .A1(F[63]), .A2(n1431), .B1(E[63]), .B2(n1425), .ZN(n29) );
  NAND4_X1 U136 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U137 ( .A1(B[41]), .A2(n1405), .B1(A[41]), .B2(n1399), .ZN(n123) );
  AOI22_X1 U138 ( .A1(D[41]), .A2(n1417), .B1(C[41]), .B2(n1411), .ZN(n124) );
  AOI22_X1 U139 ( .A1(H[41]), .A2(n1441), .B1(G[41]), .B2(n1435), .ZN(n126) );
  AOI22_X1 U140 ( .A1(D[18]), .A2(n1415), .B1(C[18]), .B2(n1409), .ZN(n228) );
  AOI22_X1 U141 ( .A1(D[17]), .A2(n1415), .B1(C[17]), .B2(n1409), .ZN(n232) );
  AOI22_X1 U142 ( .A1(D[19]), .A2(n1415), .B1(C[19]), .B2(n1409), .ZN(n224) );
  NAND4_X1 U143 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U144 ( .A1(B[39]), .A2(n1405), .B1(A[39]), .B2(n1399), .ZN(n135) );
  AOI22_X1 U145 ( .A1(D[39]), .A2(n1417), .B1(C[39]), .B2(n1411), .ZN(n136) );
  AOI22_X1 U146 ( .A1(H[39]), .A2(n1441), .B1(G[39]), .B2(n1435), .ZN(n138) );
  NAND4_X1 U147 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U148 ( .A1(B[33]), .A2(n1405), .B1(A[33]), .B2(n1399), .ZN(n159) );
  AOI22_X1 U149 ( .A1(D[33]), .A2(n1417), .B1(C[33]), .B2(n1411), .ZN(n160) );
  AOI22_X1 U150 ( .A1(H[33]), .A2(n1441), .B1(G[33]), .B2(n1435), .ZN(n162) );
  NAND4_X1 U151 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U152 ( .A1(B[28]), .A2(n1404), .B1(A[28]), .B2(n1398), .ZN(n183) );
  AOI22_X1 U153 ( .A1(D[28]), .A2(n1416), .B1(C[28]), .B2(n1410), .ZN(n184) );
  AOI22_X1 U154 ( .A1(H[28]), .A2(n1440), .B1(G[28]), .B2(n1434), .ZN(n186) );
  NAND4_X1 U155 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U156 ( .A1(H[20]), .A2(n1440), .B1(G[20]), .B2(n1434), .ZN(n218) );
  AOI22_X1 U157 ( .A1(B[20]), .A2(n1404), .B1(A[20]), .B2(n1398), .ZN(n215) );
  AOI22_X1 U158 ( .A1(D[20]), .A2(n1416), .B1(C[20]), .B2(n1410), .ZN(n216) );
  NAND4_X1 U159 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U160 ( .A1(B[22]), .A2(n1404), .B1(A[22]), .B2(n1398), .ZN(n207) );
  AOI22_X1 U161 ( .A1(H[22]), .A2(n1440), .B1(G[22]), .B2(n1434), .ZN(n210) );
  AOI22_X1 U162 ( .A1(D[22]), .A2(n1416), .B1(C[22]), .B2(n1410), .ZN(n208) );
  NAND4_X1 U163 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U164 ( .A1(H[18]), .A2(n1439), .B1(G[18]), .B2(n1433), .ZN(n230) );
  AOI22_X1 U165 ( .A1(B[18]), .A2(n1403), .B1(A[18]), .B2(n1397), .ZN(n227) );
  AOI22_X1 U166 ( .A1(F[18]), .A2(n1427), .B1(E[18]), .B2(n1421), .ZN(n229) );
  NAND4_X1 U167 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U168 ( .A1(B[31]), .A2(n1405), .B1(A[31]), .B2(n1399), .ZN(n167) );
  AOI22_X1 U169 ( .A1(D[31]), .A2(n1417), .B1(C[31]), .B2(n1411), .ZN(n168) );
  AOI22_X1 U170 ( .A1(H[31]), .A2(n1441), .B1(G[31]), .B2(n1435), .ZN(n170) );
  NAND4_X1 U171 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U172 ( .A1(B[43]), .A2(n1406), .B1(A[43]), .B2(n1400), .ZN(n115) );
  AOI22_X1 U173 ( .A1(D[43]), .A2(n1418), .B1(C[43]), .B2(n1412), .ZN(n116) );
  AOI22_X1 U174 ( .A1(H[43]), .A2(n1442), .B1(G[43]), .B2(n1436), .ZN(n118) );
  NAND4_X1 U175 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U176 ( .A1(D[16]), .A2(n1415), .B1(C[16]), .B2(n1409), .ZN(n236) );
  AOI22_X1 U177 ( .A1(H[16]), .A2(n1439), .B1(G[16]), .B2(n1433), .ZN(n238) );
  AOI22_X1 U178 ( .A1(B[16]), .A2(n1403), .B1(A[16]), .B2(n1397), .ZN(n235) );
  NAND4_X1 U179 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U180 ( .A1(B[32]), .A2(n1405), .B1(A[32]), .B2(n1399), .ZN(n163) );
  AOI22_X1 U181 ( .A1(D[32]), .A2(n1417), .B1(C[32]), .B2(n1411), .ZN(n164) );
  AOI22_X1 U182 ( .A1(H[32]), .A2(n1441), .B1(G[32]), .B2(n1435), .ZN(n166) );
  NAND4_X1 U183 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U184 ( .A1(B[38]), .A2(n1405), .B1(A[38]), .B2(n1399), .ZN(n139) );
  AOI22_X1 U185 ( .A1(D[38]), .A2(n1417), .B1(C[38]), .B2(n1411), .ZN(n140) );
  AOI22_X1 U186 ( .A1(H[38]), .A2(n1441), .B1(G[38]), .B2(n1435), .ZN(n142) );
  NAND4_X1 U187 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U188 ( .A1(B[42]), .A2(n1406), .B1(A[42]), .B2(n1400), .ZN(n119) );
  AOI22_X1 U189 ( .A1(D[42]), .A2(n1418), .B1(C[42]), .B2(n1412), .ZN(n120) );
  AOI22_X1 U190 ( .A1(H[42]), .A2(n1442), .B1(G[42]), .B2(n1436), .ZN(n122) );
  NAND4_X1 U191 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U192 ( .A1(B[45]), .A2(n1406), .B1(A[45]), .B2(n1400), .ZN(n107) );
  AOI22_X1 U193 ( .A1(D[45]), .A2(n1418), .B1(C[45]), .B2(n1412), .ZN(n108) );
  AOI22_X1 U194 ( .A1(H[45]), .A2(n1442), .B1(G[45]), .B2(n1436), .ZN(n110) );
  NAND4_X1 U195 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U196 ( .A1(B[50]), .A2(n1406), .B1(A[50]), .B2(n1400), .ZN(n83) );
  AOI22_X1 U197 ( .A1(D[50]), .A2(n1418), .B1(C[50]), .B2(n1412), .ZN(n84) );
  AOI22_X1 U198 ( .A1(H[50]), .A2(n1442), .B1(G[50]), .B2(n1436), .ZN(n86) );
  NAND4_X1 U199 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U200 ( .A1(B[48]), .A2(n1406), .B1(A[48]), .B2(n1400), .ZN(n95) );
  AOI22_X1 U201 ( .A1(D[48]), .A2(n1418), .B1(C[48]), .B2(n1412), .ZN(n96) );
  AOI22_X1 U202 ( .A1(H[48]), .A2(n1442), .B1(G[48]), .B2(n1436), .ZN(n98) );
  NAND4_X1 U203 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U204 ( .A1(B[54]), .A2(n1407), .B1(A[54]), .B2(n1401), .ZN(n67) );
  AOI22_X1 U205 ( .A1(D[54]), .A2(n1419), .B1(C[54]), .B2(n1413), .ZN(n68) );
  AOI22_X1 U206 ( .A1(H[54]), .A2(n1443), .B1(G[54]), .B2(n1437), .ZN(n70) );
  NAND4_X1 U207 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U208 ( .A1(B[58]), .A2(n1407), .B1(A[58]), .B2(n1401), .ZN(n51) );
  AOI22_X1 U209 ( .A1(D[58]), .A2(n1419), .B1(C[58]), .B2(n1413), .ZN(n52) );
  AOI22_X1 U210 ( .A1(H[58]), .A2(n1443), .B1(G[58]), .B2(n1437), .ZN(n54) );
  NAND4_X1 U211 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U212 ( .A1(B[61]), .A2(n1407), .B1(A[61]), .B2(n1401), .ZN(n35) );
  AOI22_X1 U213 ( .A1(D[61]), .A2(n1419), .B1(C[61]), .B2(n1413), .ZN(n36) );
  AOI22_X1 U214 ( .A1(H[61]), .A2(n1443), .B1(G[61]), .B2(n1437), .ZN(n38) );
  NAND4_X1 U215 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U216 ( .A1(B[63]), .A2(n1407), .B1(A[63]), .B2(n1401), .ZN(n27) );
  AOI22_X1 U217 ( .A1(D[63]), .A2(n1419), .B1(C[63]), .B2(n1413), .ZN(n28) );
  AOI22_X1 U218 ( .A1(H[63]), .A2(n1443), .B1(G[63]), .B2(n1437), .ZN(n30) );
  NAND4_X1 U219 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U220 ( .A1(B[62]), .A2(n1407), .B1(A[62]), .B2(n1401), .ZN(n31) );
  AOI22_X1 U221 ( .A1(D[62]), .A2(n1419), .B1(C[62]), .B2(n1413), .ZN(n32) );
  AOI22_X1 U222 ( .A1(H[62]), .A2(n1443), .B1(G[62]), .B2(n1437), .ZN(n34) );
  NAND4_X1 U223 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U224 ( .A1(B[25]), .A2(n1404), .B1(A[25]), .B2(n1398), .ZN(n195) );
  AOI22_X1 U225 ( .A1(D[25]), .A2(n1416), .B1(C[25]), .B2(n1410), .ZN(n196) );
  AOI22_X1 U226 ( .A1(H[25]), .A2(n1440), .B1(G[25]), .B2(n1434), .ZN(n198) );
  NAND4_X1 U227 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U228 ( .A1(B[21]), .A2(n1404), .B1(A[21]), .B2(n1398), .ZN(n211) );
  AOI22_X1 U229 ( .A1(H[21]), .A2(n1440), .B1(G[21]), .B2(n1434), .ZN(n214) );
  AOI22_X1 U230 ( .A1(D[21]), .A2(n1416), .B1(C[21]), .B2(n1410), .ZN(n212) );
  NAND4_X1 U231 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U232 ( .A1(B[29]), .A2(n1404), .B1(A[29]), .B2(n1398), .ZN(n179) );
  AOI22_X1 U233 ( .A1(D[29]), .A2(n1416), .B1(C[29]), .B2(n1410), .ZN(n180) );
  AOI22_X1 U234 ( .A1(H[29]), .A2(n1440), .B1(G[29]), .B2(n1434), .ZN(n182) );
  AOI22_X1 U235 ( .A1(F[40]), .A2(n1429), .B1(E[40]), .B2(n1423), .ZN(n129) );
  AOI22_X1 U236 ( .A1(F[44]), .A2(n1430), .B1(E[44]), .B2(n1424), .ZN(n113) );
  AOI22_X1 U237 ( .A1(F[60]), .A2(n1431), .B1(E[60]), .B2(n1425), .ZN(n41) );
  AOI22_X1 U238 ( .A1(F[58]), .A2(n1431), .B1(E[58]), .B2(n1425), .ZN(n53) );
  NAND4_X1 U239 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U240 ( .A1(B[30]), .A2(n1404), .B1(A[30]), .B2(n1398), .ZN(n171) );
  AOI22_X1 U241 ( .A1(D[30]), .A2(n1416), .B1(C[30]), .B2(n1410), .ZN(n172) );
  AOI22_X1 U242 ( .A1(H[30]), .A2(n1440), .B1(G[30]), .B2(n1434), .ZN(n174) );
  NAND4_X1 U243 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U244 ( .A1(B[36]), .A2(n1405), .B1(A[36]), .B2(n1399), .ZN(n147) );
  AOI22_X1 U245 ( .A1(D[36]), .A2(n1417), .B1(C[36]), .B2(n1411), .ZN(n148) );
  AOI22_X1 U246 ( .A1(H[36]), .A2(n1441), .B1(G[36]), .B2(n1435), .ZN(n150) );
  NAND4_X1 U247 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U248 ( .A1(B[49]), .A2(n1406), .B1(A[49]), .B2(n1400), .ZN(n91) );
  AOI22_X1 U249 ( .A1(D[49]), .A2(n1418), .B1(C[49]), .B2(n1412), .ZN(n92) );
  AOI22_X1 U250 ( .A1(H[49]), .A2(n1442), .B1(G[49]), .B2(n1436), .ZN(n94) );
  NAND4_X1 U251 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U252 ( .A1(B[51]), .A2(n1406), .B1(A[51]), .B2(n1400), .ZN(n79) );
  AOI22_X1 U253 ( .A1(D[51]), .A2(n1418), .B1(C[51]), .B2(n1412), .ZN(n80) );
  AOI22_X1 U254 ( .A1(H[51]), .A2(n1442), .B1(G[51]), .B2(n1436), .ZN(n82) );
  NAND4_X1 U255 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U256 ( .A1(B[53]), .A2(n1407), .B1(A[53]), .B2(n1401), .ZN(n71) );
  AOI22_X1 U257 ( .A1(D[53]), .A2(n1419), .B1(C[53]), .B2(n1413), .ZN(n72) );
  AOI22_X1 U258 ( .A1(H[53]), .A2(n1443), .B1(G[53]), .B2(n1437), .ZN(n74) );
  NAND4_X1 U259 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U260 ( .A1(B[52]), .A2(n1406), .B1(A[52]), .B2(n1400), .ZN(n75) );
  AOI22_X1 U261 ( .A1(D[52]), .A2(n1418), .B1(C[52]), .B2(n1412), .ZN(n76) );
  AOI22_X1 U262 ( .A1(H[52]), .A2(n1442), .B1(G[52]), .B2(n1436), .ZN(n78) );
  NAND4_X1 U263 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U264 ( .A1(B[56]), .A2(n1407), .B1(A[56]), .B2(n1401), .ZN(n59) );
  AOI22_X1 U265 ( .A1(D[56]), .A2(n1419), .B1(C[56]), .B2(n1413), .ZN(n60) );
  AOI22_X1 U266 ( .A1(H[56]), .A2(n1443), .B1(G[56]), .B2(n1437), .ZN(n62) );
  NAND4_X1 U267 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U268 ( .A1(B[57]), .A2(n1407), .B1(A[57]), .B2(n1401), .ZN(n55) );
  AOI22_X1 U269 ( .A1(D[57]), .A2(n1419), .B1(C[57]), .B2(n1413), .ZN(n56) );
  AOI22_X1 U270 ( .A1(H[57]), .A2(n1443), .B1(G[57]), .B2(n1437), .ZN(n58) );
  NAND4_X1 U271 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U272 ( .A1(H[17]), .A2(n1439), .B1(G[17]), .B2(n1433), .ZN(n234) );
  AOI22_X1 U273 ( .A1(B[17]), .A2(n1403), .B1(A[17]), .B2(n1397), .ZN(n231) );
  AOI22_X1 U274 ( .A1(F[17]), .A2(n1427), .B1(E[17]), .B2(n1421), .ZN(n233) );
  NAND4_X1 U275 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U276 ( .A1(B[44]), .A2(n1406), .B1(A[44]), .B2(n1400), .ZN(n111) );
  AOI22_X1 U277 ( .A1(D[44]), .A2(n1418), .B1(C[44]), .B2(n1412), .ZN(n112) );
  AOI22_X1 U278 ( .A1(H[44]), .A2(n1442), .B1(G[44]), .B2(n1436), .ZN(n114) );
  NAND4_X1 U279 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U280 ( .A1(B[59]), .A2(n1407), .B1(A[59]), .B2(n1401), .ZN(n47) );
  AOI22_X1 U281 ( .A1(D[59]), .A2(n1419), .B1(C[59]), .B2(n1413), .ZN(n48) );
  AOI22_X1 U282 ( .A1(H[59]), .A2(n1443), .B1(G[59]), .B2(n1437), .ZN(n50) );
  NAND4_X1 U283 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U284 ( .A1(B[60]), .A2(n1407), .B1(A[60]), .B2(n1401), .ZN(n39) );
  AOI22_X1 U285 ( .A1(D[60]), .A2(n1419), .B1(C[60]), .B2(n1413), .ZN(n40) );
  AOI22_X1 U286 ( .A1(H[60]), .A2(n1443), .B1(G[60]), .B2(n1437), .ZN(n42) );
  NAND4_X1 U287 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U288 ( .A1(B[55]), .A2(n1407), .B1(A[55]), .B2(n1401), .ZN(n63) );
  AOI22_X1 U289 ( .A1(D[55]), .A2(n1419), .B1(C[55]), .B2(n1413), .ZN(n64) );
  AOI22_X1 U290 ( .A1(H[55]), .A2(n1443), .B1(G[55]), .B2(n1437), .ZN(n66) );
  NAND4_X1 U291 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U292 ( .A1(B[0]), .A2(n1403), .B1(A[0]), .B2(n1397), .ZN(n263) );
  AOI22_X1 U293 ( .A1(D[0]), .A2(n1415), .B1(C[0]), .B2(n1409), .ZN(n264) );
  AOI22_X1 U294 ( .A1(F[0]), .A2(n1427), .B1(E[0]), .B2(n1421), .ZN(n265) );
  AOI22_X1 U295 ( .A1(H[5]), .A2(n1443), .B1(G[5]), .B2(n1437), .ZN(n46) );
  AOI22_X1 U296 ( .A1(H[13]), .A2(n1439), .B1(G[13]), .B2(n1433), .ZN(n250) );
  AOI22_X1 U297 ( .A1(H[9]), .A2(n1444), .B1(G[9]), .B2(n1438), .ZN(n6) );
  AOI22_X1 U298 ( .A1(H[7]), .A2(n1444), .B1(G[7]), .B2(n1438), .ZN(n22) );
  AOI22_X1 U299 ( .A1(H[11]), .A2(n1439), .B1(G[11]), .B2(n1433), .ZN(n258) );
  AOI22_X1 U300 ( .A1(H[15]), .A2(n1439), .B1(G[15]), .B2(n1433), .ZN(n242) );
  AOI22_X1 U301 ( .A1(H[3]), .A2(n1441), .B1(G[3]), .B2(n1435), .ZN(n134) );
  AOI22_X1 U302 ( .A1(H[4]), .A2(n1442), .B1(G[4]), .B2(n1436), .ZN(n90) );
  AOI22_X1 U303 ( .A1(H[12]), .A2(n1439), .B1(G[12]), .B2(n1433), .ZN(n254) );
  AOI22_X1 U304 ( .A1(H[8]), .A2(n1444), .B1(G[8]), .B2(n1438), .ZN(n18) );
  AOI22_X1 U305 ( .A1(H[6]), .A2(n1444), .B1(G[6]), .B2(n1438), .ZN(n26) );
  AOI22_X1 U306 ( .A1(H[10]), .A2(n1439), .B1(G[10]), .B2(n1433), .ZN(n262) );
  AOI22_X1 U307 ( .A1(H[14]), .A2(n1439), .B1(G[14]), .B2(n1433), .ZN(n246) );
  AOI22_X1 U308 ( .A1(H[2]), .A2(n1440), .B1(G[2]), .B2(n1434), .ZN(n178) );
  AOI22_X1 U309 ( .A1(H[1]), .A2(n1439), .B1(G[1]), .B2(n1433), .ZN(n222) );
  NAND4_X1 U310 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U311 ( .A1(B[4]), .A2(n1406), .B1(A[4]), .B2(n1400), .ZN(n87) );
  AOI22_X1 U312 ( .A1(D[4]), .A2(n1418), .B1(C[4]), .B2(n1412), .ZN(n88) );
  AOI22_X1 U313 ( .A1(F[4]), .A2(n1430), .B1(E[4]), .B2(n1424), .ZN(n89) );
  NAND4_X1 U314 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U315 ( .A1(B[5]), .A2(n1407), .B1(A[5]), .B2(n1401), .ZN(n43) );
  AOI22_X1 U316 ( .A1(D[5]), .A2(n1419), .B1(C[5]), .B2(n1413), .ZN(n44) );
  AOI22_X1 U317 ( .A1(F[5]), .A2(n1431), .B1(E[5]), .B2(n1425), .ZN(n45) );
  NAND4_X1 U318 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U319 ( .A1(B[12]), .A2(n1403), .B1(A[12]), .B2(n1397), .ZN(n251) );
  AOI22_X1 U320 ( .A1(D[12]), .A2(n1415), .B1(C[12]), .B2(n1409), .ZN(n252) );
  AOI22_X1 U321 ( .A1(F[12]), .A2(n1427), .B1(E[12]), .B2(n1421), .ZN(n253) );
  NAND4_X1 U322 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U323 ( .A1(B[13]), .A2(n1403), .B1(A[13]), .B2(n1397), .ZN(n247) );
  AOI22_X1 U324 ( .A1(D[13]), .A2(n1415), .B1(C[13]), .B2(n1409), .ZN(n248) );
  AOI22_X1 U325 ( .A1(F[13]), .A2(n1427), .B1(E[13]), .B2(n1421), .ZN(n249) );
  NAND4_X1 U326 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U327 ( .A1(B[8]), .A2(n1408), .B1(A[8]), .B2(n1402), .ZN(n15) );
  AOI22_X1 U328 ( .A1(D[8]), .A2(n1420), .B1(C[8]), .B2(n1414), .ZN(n16) );
  AOI22_X1 U329 ( .A1(F[8]), .A2(n1432), .B1(E[8]), .B2(n1426), .ZN(n17) );
  NAND4_X1 U330 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U331 ( .A1(B[9]), .A2(n1408), .B1(A[9]), .B2(n1402), .ZN(n3) );
  AOI22_X1 U332 ( .A1(D[9]), .A2(n1420), .B1(C[9]), .B2(n1414), .ZN(n4) );
  AOI22_X1 U333 ( .A1(F[9]), .A2(n1432), .B1(E[9]), .B2(n1426), .ZN(n5) );
  NAND4_X1 U334 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U335 ( .A1(B[11]), .A2(n1403), .B1(A[11]), .B2(n1397), .ZN(n255) );
  AOI22_X1 U336 ( .A1(D[11]), .A2(n1415), .B1(C[11]), .B2(n1409), .ZN(n256) );
  AOI22_X1 U337 ( .A1(F[11]), .A2(n1427), .B1(E[11]), .B2(n1421), .ZN(n257) );
  NAND4_X1 U338 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U339 ( .A1(B[15]), .A2(n1403), .B1(A[15]), .B2(n1397), .ZN(n239) );
  AOI22_X1 U340 ( .A1(D[15]), .A2(n1415), .B1(C[15]), .B2(n1409), .ZN(n240) );
  AOI22_X1 U341 ( .A1(F[15]), .A2(n1427), .B1(E[15]), .B2(n1421), .ZN(n241) );
  NAND4_X1 U342 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U343 ( .A1(B[7]), .A2(n1408), .B1(A[7]), .B2(n1402), .ZN(n19) );
  AOI22_X1 U344 ( .A1(D[7]), .A2(n1420), .B1(C[7]), .B2(n1414), .ZN(n20) );
  AOI22_X1 U345 ( .A1(F[7]), .A2(n1432), .B1(E[7]), .B2(n1426), .ZN(n21) );
  NAND4_X1 U346 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U347 ( .A1(B[6]), .A2(n1408), .B1(A[6]), .B2(n1402), .ZN(n23) );
  AOI22_X1 U348 ( .A1(D[6]), .A2(n1420), .B1(C[6]), .B2(n1414), .ZN(n24) );
  AOI22_X1 U349 ( .A1(F[6]), .A2(n1432), .B1(E[6]), .B2(n1426), .ZN(n25) );
  NAND4_X1 U350 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U351 ( .A1(B[10]), .A2(n1403), .B1(A[10]), .B2(n1397), .ZN(n259) );
  AOI22_X1 U352 ( .A1(D[10]), .A2(n1415), .B1(C[10]), .B2(n1409), .ZN(n260) );
  AOI22_X1 U353 ( .A1(F[10]), .A2(n1427), .B1(E[10]), .B2(n1421), .ZN(n261) );
  NAND4_X1 U354 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U355 ( .A1(B[14]), .A2(n1403), .B1(A[14]), .B2(n1397), .ZN(n243) );
  AOI22_X1 U356 ( .A1(D[14]), .A2(n1415), .B1(C[14]), .B2(n1409), .ZN(n244) );
  AOI22_X1 U357 ( .A1(F[14]), .A2(n1427), .B1(E[14]), .B2(n1421), .ZN(n245) );
  NAND4_X1 U358 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U359 ( .A1(B[3]), .A2(n1405), .B1(A[3]), .B2(n1399), .ZN(n131) );
  AOI22_X1 U360 ( .A1(D[3]), .A2(n1417), .B1(C[3]), .B2(n1411), .ZN(n132) );
  AOI22_X1 U361 ( .A1(F[3]), .A2(n1429), .B1(E[3]), .B2(n1423), .ZN(n133) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1404), .B1(A[2]), .B2(n1398), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1416), .B1(C[2]), .B2(n1410), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1428), .B1(E[2]), .B2(n1422), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1403), .B1(A[1]), .B2(n1397), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1415), .B1(C[1]), .B2(n1409), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1427), .B1(E[1]), .B2(n1421), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1439), .B1(G[0]), .B2(n1433), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1402) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1408) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1414) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1420) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1426) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1432) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1438) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1444) );
endmodule


module MUX81_GENERIC_NBIT64_7 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n13), .Z(n1408) );
  BUF_X1 U2 ( .A(n13), .Z(n1407) );
  BUF_X1 U3 ( .A(n12), .Z(n1414) );
  BUF_X1 U4 ( .A(n12), .Z(n1413) );
  BUF_X1 U5 ( .A(n8), .Z(n1438) );
  BUF_X1 U6 ( .A(n8), .Z(n1437) );
  BUF_X1 U7 ( .A(n10), .Z(n1426) );
  BUF_X1 U8 ( .A(n10), .Z(n1425) );
  BUF_X1 U9 ( .A(n13), .Z(n1410) );
  BUF_X1 U10 ( .A(n13), .Z(n1409) );
  BUF_X1 U11 ( .A(n12), .Z(n1416) );
  BUF_X1 U12 ( .A(n12), .Z(n1415) );
  BUF_X1 U13 ( .A(n8), .Z(n1439) );
  BUF_X1 U14 ( .A(n10), .Z(n1428) );
  BUF_X1 U15 ( .A(n8), .Z(n1440) );
  BUF_X1 U16 ( .A(n10), .Z(n1427) );
  BUF_X1 U17 ( .A(n13), .Z(n1411) );
  BUF_X1 U18 ( .A(n12), .Z(n1417) );
  BUF_X1 U19 ( .A(n10), .Z(n1429) );
  BUF_X1 U20 ( .A(n8), .Z(n1441) );
  BUF_X1 U21 ( .A(n11), .Z(n1422) );
  BUF_X1 U22 ( .A(n11), .Z(n1423) );
  BUF_X1 U23 ( .A(n11), .Z(n1420) );
  BUF_X1 U24 ( .A(n11), .Z(n1421) );
  BUF_X1 U25 ( .A(n11), .Z(n1419) );
  BUF_X1 U26 ( .A(n7), .Z(n1444) );
  BUF_X1 U27 ( .A(n7), .Z(n1445) );
  BUF_X1 U28 ( .A(n9), .Z(n1434) );
  BUF_X1 U29 ( .A(n7), .Z(n1446) );
  BUF_X1 U30 ( .A(n7), .Z(n1443) );
  BUF_X1 U31 ( .A(n9), .Z(n1435) );
  BUF_X1 U32 ( .A(n7), .Z(n1447) );
  BUF_X1 U33 ( .A(n9), .Z(n1432) );
  BUF_X1 U34 ( .A(n9), .Z(n1433) );
  BUF_X1 U35 ( .A(n9), .Z(n1431) );
  BUF_X1 U36 ( .A(n14), .Z(n1404) );
  BUF_X1 U37 ( .A(n14), .Z(n1405) );
  BUF_X1 U38 ( .A(n14), .Z(n1402) );
  BUF_X1 U39 ( .A(n14), .Z(n1403) );
  BUF_X1 U40 ( .A(n14), .Z(n1401) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1449) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U52 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U53 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U54 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  NAND4_X1 U55 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U56 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U57 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U58 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  AOI22_X1 U59 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  AOI22_X1 U60 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  AOI22_X1 U61 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  AOI22_X1 U62 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U63 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U64 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  NAND4_X1 U65 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U66 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U67 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  AOI22_X1 U68 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  NAND4_X1 U69 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U70 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U71 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  AOI22_X1 U72 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  NAND4_X1 U73 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U74 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U75 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U76 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  NAND4_X1 U77 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U78 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U79 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U80 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  NAND4_X1 U81 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U82 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U83 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U84 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  NAND4_X1 U85 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U86 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U87 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U88 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  NAND4_X1 U89 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U90 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U91 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U92 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  NAND4_X1 U93 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U94 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U95 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U96 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  NAND4_X1 U97 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U98 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U99 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U100 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  AOI22_X1 U101 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  AOI22_X1 U102 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  AOI22_X1 U103 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  AOI22_X1 U104 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  AOI22_X1 U105 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  AOI22_X1 U106 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  AOI22_X1 U107 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  AOI22_X1 U108 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  AOI22_X1 U109 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  AOI22_X1 U110 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  AOI22_X1 U111 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  AOI22_X1 U112 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  AOI22_X1 U113 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  AOI22_X1 U114 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  AOI22_X1 U115 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  AOI22_X1 U116 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  AOI22_X1 U117 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  AOI22_X1 U118 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  AOI22_X1 U119 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  AOI22_X1 U120 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  AOI22_X1 U121 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  AOI22_X1 U122 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  AOI22_X1 U123 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  AOI22_X1 U124 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  AOI22_X1 U125 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  AOI22_X1 U126 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  AOI22_X1 U127 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  AOI22_X1 U128 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  AOI22_X1 U129 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  AOI22_X1 U130 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  AOI22_X1 U131 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U132 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U133 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U134 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U135 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  AOI22_X1 U136 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  AOI22_X1 U137 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  AOI22_X1 U138 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  AOI22_X1 U139 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  AOI22_X1 U140 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  AOI22_X1 U141 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  NAND4_X1 U142 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U143 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U144 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U145 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  NAND4_X1 U146 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U147 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U148 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U149 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  NAND4_X1 U150 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U151 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  AOI22_X1 U152 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U153 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  NAND4_X1 U154 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U155 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U156 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U157 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  NAND4_X1 U158 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U159 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U160 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U161 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  NAND4_X1 U162 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U163 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U164 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  AOI22_X1 U165 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  NAND4_X1 U166 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U167 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U168 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U169 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  NAND4_X1 U170 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U171 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U172 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U173 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  NAND4_X1 U174 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U175 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U176 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  AOI22_X1 U177 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  NAND4_X1 U178 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U179 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U180 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  AOI22_X1 U181 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  NAND4_X1 U182 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U183 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U184 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U185 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  NAND4_X1 U186 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U187 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U188 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U189 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  NAND4_X1 U190 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U191 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U192 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U193 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  NAND4_X1 U194 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U195 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U196 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U197 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  NAND4_X1 U198 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U199 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U200 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U201 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  NAND4_X1 U202 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U203 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U204 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U205 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  NAND4_X1 U206 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U207 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U208 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U209 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  NAND4_X1 U210 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U211 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U212 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U213 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  NAND4_X1 U214 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U215 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U216 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U217 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  NAND4_X1 U218 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U219 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U220 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U221 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  NAND4_X1 U222 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U223 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U224 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U225 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  AOI22_X1 U226 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  NAND4_X1 U227 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U228 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U229 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U230 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  NAND4_X1 U231 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U232 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U233 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U234 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  AOI22_X1 U235 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  AOI22_X1 U236 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  AOI22_X1 U237 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  NAND4_X1 U238 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U239 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U240 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  AOI22_X1 U241 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  NAND4_X1 U242 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U243 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U244 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U245 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  NAND4_X1 U246 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U247 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U248 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U249 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  NAND4_X1 U250 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U251 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U252 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U253 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  NAND4_X1 U254 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U255 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  AOI22_X1 U256 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  AOI22_X1 U257 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  NAND4_X1 U258 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U259 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U260 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U261 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  NAND4_X1 U262 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U263 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U264 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U265 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  NAND4_X1 U266 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U267 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U268 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U269 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  NAND4_X1 U270 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U271 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  AOI22_X1 U272 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U273 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  AOI22_X1 U274 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  AOI22_X1 U275 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  NAND4_X1 U276 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U277 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U278 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U279 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  NAND4_X1 U280 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U281 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U282 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U283 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U284 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U285 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U286 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U287 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U288 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U289 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U290 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  AOI22_X1 U291 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U292 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U293 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U294 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U295 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U296 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U297 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U298 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U299 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U300 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U301 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U302 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U303 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U304 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U305 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U306 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U307 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U308 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U309 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U310 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U311 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U312 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U313 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U314 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U315 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U316 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U317 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U318 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U319 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  AOI22_X1 U320 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  NAND4_X1 U321 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U322 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U323 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U324 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U325 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U326 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  AOI22_X1 U327 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  AOI22_X1 U328 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  NAND4_X1 U329 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U330 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U331 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  AOI22_X1 U332 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  NAND4_X1 U333 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U334 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U335 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U336 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U337 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U338 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U339 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U340 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U341 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U342 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U343 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  AOI22_X1 U344 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  NAND4_X1 U345 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U346 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U347 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U348 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U349 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U350 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U351 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U352 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U353 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U354 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  AOI22_X1 U355 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  AOI22_X1 U356 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  NAND4_X1 U357 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U358 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U359 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U360 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U361 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U362 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U363 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U364 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U365 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U366 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U367 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U368 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U369 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  NAND4_X1 U370 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_6 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n13), .Z(n1408) );
  BUF_X1 U2 ( .A(n13), .Z(n1409) );
  BUF_X1 U3 ( .A(n12), .Z(n1416) );
  BUF_X1 U4 ( .A(n12), .Z(n1414) );
  BUF_X1 U5 ( .A(n12), .Z(n1415) );
  BUF_X1 U6 ( .A(n8), .Z(n1438) );
  BUF_X1 U7 ( .A(n8), .Z(n1439) );
  BUF_X1 U8 ( .A(n10), .Z(n1428) );
  BUF_X1 U9 ( .A(n10), .Z(n1426) );
  BUF_X1 U10 ( .A(n10), .Z(n1427) );
  BUF_X1 U11 ( .A(n13), .Z(n1410) );
  BUF_X1 U12 ( .A(n13), .Z(n1411) );
  BUF_X1 U13 ( .A(n12), .Z(n1417) );
  BUF_X1 U14 ( .A(n8), .Z(n1440) );
  BUF_X1 U15 ( .A(n10), .Z(n1429) );
  BUF_X1 U16 ( .A(n8), .Z(n1441) );
  BUF_X1 U17 ( .A(n11), .Z(n1422) );
  BUF_X1 U18 ( .A(n11), .Z(n1420) );
  BUF_X1 U19 ( .A(n11), .Z(n1421) );
  BUF_X1 U20 ( .A(n11), .Z(n1419) );
  BUF_X1 U21 ( .A(n13), .Z(n1407) );
  BUF_X1 U22 ( .A(n11), .Z(n1423) );
  BUF_X1 U23 ( .A(n7), .Z(n1443) );
  BUF_X1 U24 ( .A(n7), .Z(n1444) );
  BUF_X1 U25 ( .A(n7), .Z(n1445) );
  BUF_X1 U26 ( .A(n9), .Z(n1434) );
  BUF_X1 U27 ( .A(n7), .Z(n1446) );
  BUF_X1 U28 ( .A(n9), .Z(n1435) );
  BUF_X1 U29 ( .A(n9), .Z(n1432) );
  BUF_X1 U30 ( .A(n9), .Z(n1433) );
  BUF_X1 U31 ( .A(n9), .Z(n1431) );
  BUF_X1 U32 ( .A(n7), .Z(n1447) );
  BUF_X1 U33 ( .A(n14), .Z(n1404) );
  BUF_X1 U34 ( .A(n14), .Z(n1402) );
  BUF_X1 U35 ( .A(n14), .Z(n1403) );
  BUF_X1 U36 ( .A(n12), .Z(n1413) );
  BUF_X1 U37 ( .A(n14), .Z(n1401) );
  BUF_X1 U38 ( .A(n14), .Z(n1405) );
  BUF_X1 U39 ( .A(n8), .Z(n1437) );
  BUF_X1 U40 ( .A(n10), .Z(n1425) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1449) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  AOI22_X1 U51 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  AOI22_X1 U52 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  AOI22_X1 U53 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  NAND4_X1 U54 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U55 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U56 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U57 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  NAND4_X1 U58 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U59 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U60 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U61 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  NAND4_X1 U62 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U63 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U64 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U65 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  NAND4_X1 U66 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U67 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U68 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U69 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  AOI22_X1 U70 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  AOI22_X1 U71 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  AOI22_X1 U72 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  AOI22_X1 U73 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  AOI22_X1 U74 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  AOI22_X1 U75 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  AOI22_X1 U76 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  AOI22_X1 U77 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  AOI22_X1 U78 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  AOI22_X1 U79 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  AOI22_X1 U80 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  AOI22_X1 U81 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  AOI22_X1 U82 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  AOI22_X1 U83 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  AOI22_X1 U84 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  AOI22_X1 U85 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  AOI22_X1 U86 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  AOI22_X1 U87 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  AOI22_X1 U88 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  AOI22_X1 U89 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U90 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U91 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U92 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U93 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  NAND4_X1 U94 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U95 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U96 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U97 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  NAND4_X1 U98 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U99 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U100 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U101 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  NAND4_X1 U102 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U103 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U104 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U105 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  NAND4_X1 U106 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U107 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U108 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U109 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  NAND4_X1 U110 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U111 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U112 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U113 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  NAND4_X1 U114 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U115 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U116 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U117 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  NAND4_X1 U118 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U119 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U120 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U121 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  NAND4_X1 U122 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U123 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U124 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U125 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  NAND4_X1 U126 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U127 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U128 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U129 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  NAND4_X1 U130 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U131 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U132 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U133 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  AOI22_X1 U134 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  NAND4_X1 U135 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U136 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U137 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U138 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  AOI22_X1 U139 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  AOI22_X1 U140 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  NAND4_X1 U141 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U142 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U143 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U144 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  NAND4_X1 U145 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U146 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U147 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U148 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  NAND4_X1 U149 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U150 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U151 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U152 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  NAND4_X1 U153 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U154 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U155 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U156 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  NAND4_X1 U157 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U158 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U159 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U160 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  NAND4_X1 U161 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U162 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U163 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U164 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  NAND4_X1 U165 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U166 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U167 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U168 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  NAND4_X1 U169 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U170 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U171 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U172 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  NAND4_X1 U173 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U174 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U175 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U176 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  NAND4_X1 U177 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U178 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U179 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U180 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  NAND4_X1 U181 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U182 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U183 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U184 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  NAND4_X1 U185 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U186 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U187 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U188 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  NAND4_X1 U189 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U190 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U191 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U192 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  AOI22_X1 U193 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  AOI22_X1 U194 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  AOI22_X1 U195 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  AOI22_X1 U196 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  AOI22_X1 U197 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  AOI22_X1 U198 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  AOI22_X1 U199 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  AOI22_X1 U200 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  AOI22_X1 U201 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  AOI22_X1 U202 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  AOI22_X1 U203 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  AOI22_X1 U204 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  AOI22_X1 U205 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  AOI22_X1 U206 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  NAND4_X1 U207 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U208 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U209 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  AOI22_X1 U210 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  AOI22_X1 U211 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  AOI22_X1 U212 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  AOI22_X1 U213 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  AOI22_X1 U214 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  NAND4_X1 U215 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U216 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U217 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U218 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  NAND4_X1 U219 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U220 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U221 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U222 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  NAND4_X1 U223 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U224 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U225 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U226 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  NAND4_X1 U227 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U228 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U229 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  AOI22_X1 U230 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  NAND4_X1 U231 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U232 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  AOI22_X1 U233 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U234 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  NAND4_X1 U235 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U236 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U237 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U238 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  NAND4_X1 U239 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U240 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U241 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  AOI22_X1 U242 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  NAND4_X1 U243 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U244 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U245 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  AOI22_X1 U246 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  NAND4_X1 U247 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U248 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U249 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U250 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  NAND4_X1 U251 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U252 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U253 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U254 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  NAND4_X1 U255 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U256 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U257 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U258 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  NAND4_X1 U259 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U260 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U261 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U262 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  NAND4_X1 U263 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U264 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  AOI22_X1 U265 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U266 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  NAND4_X1 U267 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U268 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U269 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  AOI22_X1 U270 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  NAND4_X1 U271 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U272 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U273 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U274 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U275 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U276 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U277 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U278 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U279 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U280 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U281 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  AOI22_X1 U282 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  AOI22_X1 U283 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U284 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U285 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U286 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U287 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U288 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U289 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U290 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U291 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  AOI22_X1 U292 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U293 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U294 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U295 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U296 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U297 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U298 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U299 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U300 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U301 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U302 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U303 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  AOI22_X1 U304 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  AOI22_X1 U305 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  NAND4_X1 U306 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U307 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U308 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  AOI22_X1 U309 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  NAND4_X1 U310 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U311 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U312 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  AOI22_X1 U313 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  NAND4_X1 U314 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U315 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U316 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U317 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U318 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U319 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U320 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U321 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U322 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U323 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U324 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U325 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U326 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U327 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U328 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U329 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U330 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U331 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U332 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  AOI22_X1 U333 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  NAND4_X1 U334 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U335 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U336 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U337 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U338 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U339 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U340 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U341 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U342 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U343 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U344 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U345 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U346 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U347 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U348 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U349 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U350 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U351 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U352 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  AOI22_X1 U353 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  NAND4_X1 U354 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U355 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  AOI22_X1 U356 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  AOI22_X1 U357 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  NAND4_X1 U358 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U359 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  AOI22_X1 U360 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  AOI22_X1 U361 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_5 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450;

  BUF_X1 U1 ( .A(n13), .Z(n1408) );
  BUF_X1 U2 ( .A(n13), .Z(n1409) );
  BUF_X1 U3 ( .A(n12), .Z(n1414) );
  BUF_X1 U4 ( .A(n12), .Z(n1415) );
  BUF_X1 U5 ( .A(n8), .Z(n1439) );
  BUF_X1 U6 ( .A(n8), .Z(n1438) );
  BUF_X1 U7 ( .A(n10), .Z(n1426) );
  BUF_X1 U8 ( .A(n10), .Z(n1427) );
  BUF_X1 U9 ( .A(n13), .Z(n1410) );
  BUF_X1 U10 ( .A(n13), .Z(n1411) );
  BUF_X1 U11 ( .A(n12), .Z(n1416) );
  BUF_X1 U12 ( .A(n12), .Z(n1417) );
  BUF_X1 U13 ( .A(n10), .Z(n1428) );
  BUF_X1 U14 ( .A(n8), .Z(n1440) );
  BUF_X1 U15 ( .A(n10), .Z(n1429) );
  BUF_X1 U16 ( .A(n8), .Z(n1441) );
  BUF_X1 U17 ( .A(n11), .Z(n1422) );
  BUF_X1 U18 ( .A(n11), .Z(n1420) );
  BUF_X1 U19 ( .A(n11), .Z(n1421) );
  BUF_X1 U20 ( .A(n11), .Z(n1419) );
  BUF_X1 U21 ( .A(n13), .Z(n1407) );
  BUF_X1 U22 ( .A(n11), .Z(n1423) );
  BUF_X1 U23 ( .A(n7), .Z(n1443) );
  BUF_X1 U24 ( .A(n7), .Z(n1445) );
  BUF_X1 U25 ( .A(n9), .Z(n1434) );
  BUF_X1 U26 ( .A(n7), .Z(n1446) );
  BUF_X1 U27 ( .A(n7), .Z(n1444) );
  BUF_X1 U28 ( .A(n9), .Z(n1435) );
  BUF_X1 U29 ( .A(n9), .Z(n1432) );
  BUF_X1 U30 ( .A(n9), .Z(n1433) );
  BUF_X1 U31 ( .A(n9), .Z(n1431) );
  BUF_X1 U32 ( .A(n7), .Z(n1447) );
  BUF_X1 U33 ( .A(n14), .Z(n1404) );
  BUF_X1 U34 ( .A(n14), .Z(n1402) );
  BUF_X1 U35 ( .A(n14), .Z(n1403) );
  BUF_X1 U36 ( .A(n12), .Z(n1413) );
  BUF_X1 U37 ( .A(n14), .Z(n1401) );
  BUF_X1 U38 ( .A(n14), .Z(n1405) );
  BUF_X1 U39 ( .A(n8), .Z(n1437) );
  BUF_X1 U40 ( .A(n10), .Z(n1425) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1449), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1450), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1450), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1450), .A2(n1449), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1449) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1450) );
  NOR3_X1 U47 ( .A1(n1450), .A2(SEL[2]), .A3(n1449), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1449), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U52 ( .A1(B[43]), .A2(n1410), .B1(A[43]), .B2(n1404), .ZN(n115) );
  AOI22_X1 U53 ( .A1(D[43]), .A2(n1422), .B1(C[43]), .B2(n1416), .ZN(n116) );
  AOI22_X1 U54 ( .A1(H[43]), .A2(n1446), .B1(G[43]), .B2(n1440), .ZN(n118) );
  NAND4_X1 U55 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U56 ( .A1(B[48]), .A2(n1410), .B1(A[48]), .B2(n1404), .ZN(n95) );
  AOI22_X1 U57 ( .A1(D[48]), .A2(n1422), .B1(C[48]), .B2(n1416), .ZN(n96) );
  AOI22_X1 U58 ( .A1(H[48]), .A2(n1446), .B1(G[48]), .B2(n1440), .ZN(n98) );
  NAND4_X1 U59 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U60 ( .A1(B[45]), .A2(n1410), .B1(A[45]), .B2(n1404), .ZN(n107) );
  AOI22_X1 U61 ( .A1(D[45]), .A2(n1422), .B1(C[45]), .B2(n1416), .ZN(n108) );
  AOI22_X1 U62 ( .A1(H[45]), .A2(n1446), .B1(G[45]), .B2(n1440), .ZN(n110) );
  AOI22_X1 U63 ( .A1(F[53]), .A2(n1435), .B1(E[53]), .B2(n1429), .ZN(n73) );
  AOI22_X1 U64 ( .A1(F[57]), .A2(n1435), .B1(E[57]), .B2(n1429), .ZN(n57) );
  AOI22_X1 U65 ( .A1(F[59]), .A2(n1435), .B1(E[59]), .B2(n1429), .ZN(n49) );
  AOI22_X1 U66 ( .A1(F[62]), .A2(n1435), .B1(E[62]), .B2(n1429), .ZN(n33) );
  AOI22_X1 U67 ( .A1(F[51]), .A2(n1434), .B1(E[51]), .B2(n1428), .ZN(n81) );
  AOI22_X1 U68 ( .A1(F[61]), .A2(n1435), .B1(E[61]), .B2(n1429), .ZN(n37) );
  NAND4_X1 U69 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U70 ( .A1(B[47]), .A2(n1410), .B1(A[47]), .B2(n1404), .ZN(n99) );
  AOI22_X1 U71 ( .A1(D[47]), .A2(n1422), .B1(C[47]), .B2(n1416), .ZN(n100) );
  AOI22_X1 U72 ( .A1(H[47]), .A2(n1446), .B1(G[47]), .B2(n1440), .ZN(n102) );
  NAND4_X1 U73 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U74 ( .A1(B[30]), .A2(n1408), .B1(A[30]), .B2(n1402), .ZN(n171) );
  AOI22_X1 U75 ( .A1(D[30]), .A2(n1420), .B1(C[30]), .B2(n1414), .ZN(n172) );
  AOI22_X1 U76 ( .A1(H[30]), .A2(n1444), .B1(G[30]), .B2(n1438), .ZN(n174) );
  NAND4_X1 U77 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U78 ( .A1(B[50]), .A2(n1410), .B1(A[50]), .B2(n1404), .ZN(n83) );
  AOI22_X1 U79 ( .A1(D[50]), .A2(n1422), .B1(C[50]), .B2(n1416), .ZN(n84) );
  AOI22_X1 U80 ( .A1(H[50]), .A2(n1446), .B1(G[50]), .B2(n1440), .ZN(n86) );
  NAND4_X1 U81 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U82 ( .A1(B[49]), .A2(n1410), .B1(A[49]), .B2(n1404), .ZN(n91) );
  AOI22_X1 U83 ( .A1(D[49]), .A2(n1422), .B1(C[49]), .B2(n1416), .ZN(n92) );
  AOI22_X1 U84 ( .A1(H[49]), .A2(n1446), .B1(G[49]), .B2(n1440), .ZN(n94) );
  NAND4_X1 U85 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U86 ( .A1(B[52]), .A2(n1410), .B1(A[52]), .B2(n1404), .ZN(n75) );
  AOI22_X1 U87 ( .A1(D[52]), .A2(n1422), .B1(C[52]), .B2(n1416), .ZN(n76) );
  AOI22_X1 U88 ( .A1(H[52]), .A2(n1446), .B1(G[52]), .B2(n1440), .ZN(n78) );
  NAND4_X1 U89 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U90 ( .A1(B[42]), .A2(n1410), .B1(A[42]), .B2(n1404), .ZN(n119) );
  AOI22_X1 U91 ( .A1(D[42]), .A2(n1422), .B1(C[42]), .B2(n1416), .ZN(n120) );
  AOI22_X1 U92 ( .A1(H[42]), .A2(n1446), .B1(G[42]), .B2(n1440), .ZN(n122) );
  NAND4_X1 U93 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U94 ( .A1(B[51]), .A2(n1410), .B1(A[51]), .B2(n1404), .ZN(n79) );
  AOI22_X1 U95 ( .A1(D[51]), .A2(n1422), .B1(C[51]), .B2(n1416), .ZN(n80) );
  AOI22_X1 U96 ( .A1(H[51]), .A2(n1446), .B1(G[51]), .B2(n1440), .ZN(n82) );
  AOI22_X1 U97 ( .A1(F[29]), .A2(n1432), .B1(E[29]), .B2(n1426), .ZN(n181) );
  AOI22_X1 U98 ( .A1(F[31]), .A2(n1433), .B1(E[31]), .B2(n1427), .ZN(n169) );
  AOI22_X1 U99 ( .A1(F[30]), .A2(n1432), .B1(E[30]), .B2(n1426), .ZN(n173) );
  AOI22_X1 U100 ( .A1(F[32]), .A2(n1433), .B1(E[32]), .B2(n1427), .ZN(n165) );
  AOI22_X1 U101 ( .A1(F[35]), .A2(n1433), .B1(E[35]), .B2(n1427), .ZN(n153) );
  AOI22_X1 U102 ( .A1(F[33]), .A2(n1433), .B1(E[33]), .B2(n1427), .ZN(n161) );
  AOI22_X1 U103 ( .A1(F[36]), .A2(n1433), .B1(E[36]), .B2(n1427), .ZN(n149) );
  AOI22_X1 U104 ( .A1(F[37]), .A2(n1433), .B1(E[37]), .B2(n1427), .ZN(n145) );
  AOI22_X1 U105 ( .A1(F[38]), .A2(n1433), .B1(E[38]), .B2(n1427), .ZN(n141) );
  AOI22_X1 U106 ( .A1(F[39]), .A2(n1433), .B1(E[39]), .B2(n1427), .ZN(n137) );
  AOI22_X1 U107 ( .A1(F[41]), .A2(n1433), .B1(E[41]), .B2(n1427), .ZN(n125) );
  AOI22_X1 U108 ( .A1(F[44]), .A2(n1434), .B1(E[44]), .B2(n1428), .ZN(n113) );
  AOI22_X1 U109 ( .A1(F[42]), .A2(n1434), .B1(E[42]), .B2(n1428), .ZN(n121) );
  AOI22_X1 U110 ( .A1(F[40]), .A2(n1433), .B1(E[40]), .B2(n1427), .ZN(n129) );
  AOI22_X1 U111 ( .A1(F[47]), .A2(n1434), .B1(E[47]), .B2(n1428), .ZN(n101) );
  AOI22_X1 U112 ( .A1(F[43]), .A2(n1434), .B1(E[43]), .B2(n1428), .ZN(n117) );
  AOI22_X1 U113 ( .A1(F[49]), .A2(n1434), .B1(E[49]), .B2(n1428), .ZN(n93) );
  AOI22_X1 U114 ( .A1(F[45]), .A2(n1434), .B1(E[45]), .B2(n1428), .ZN(n109) );
  AOI22_X1 U115 ( .A1(F[50]), .A2(n1434), .B1(E[50]), .B2(n1428), .ZN(n85) );
  AOI22_X1 U116 ( .A1(F[54]), .A2(n1435), .B1(E[54]), .B2(n1429), .ZN(n69) );
  AOI22_X1 U117 ( .A1(F[22]), .A2(n1432), .B1(E[22]), .B2(n1426), .ZN(n209) );
  AOI22_X1 U118 ( .A1(F[55]), .A2(n1435), .B1(E[55]), .B2(n1429), .ZN(n65) );
  AOI22_X1 U119 ( .A1(F[23]), .A2(n1432), .B1(E[23]), .B2(n1426), .ZN(n205) );
  AOI22_X1 U120 ( .A1(F[58]), .A2(n1435), .B1(E[58]), .B2(n1429), .ZN(n53) );
  AOI22_X1 U121 ( .A1(F[63]), .A2(n1435), .B1(E[63]), .B2(n1429), .ZN(n29) );
  NAND4_X1 U122 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U123 ( .A1(B[35]), .A2(n1409), .B1(A[35]), .B2(n1403), .ZN(n151) );
  AOI22_X1 U124 ( .A1(D[35]), .A2(n1421), .B1(C[35]), .B2(n1415), .ZN(n152) );
  AOI22_X1 U125 ( .A1(H[35]), .A2(n1445), .B1(G[35]), .B2(n1439), .ZN(n154) );
  NAND4_X1 U126 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U127 ( .A1(B[53]), .A2(n1411), .B1(A[53]), .B2(n1405), .ZN(n71) );
  AOI22_X1 U128 ( .A1(D[53]), .A2(n1423), .B1(C[53]), .B2(n1417), .ZN(n72) );
  AOI22_X1 U129 ( .A1(H[53]), .A2(n1447), .B1(G[53]), .B2(n1441), .ZN(n74) );
  AOI22_X1 U130 ( .A1(D[27]), .A2(n1420), .B1(C[27]), .B2(n1414), .ZN(n188) );
  AOI22_X1 U131 ( .A1(D[24]), .A2(n1420), .B1(C[24]), .B2(n1414), .ZN(n200) );
  AOI22_X1 U132 ( .A1(D[25]), .A2(n1420), .B1(C[25]), .B2(n1414), .ZN(n196) );
  AOI22_X1 U133 ( .A1(D[28]), .A2(n1420), .B1(C[28]), .B2(n1414), .ZN(n184) );
  AOI22_X1 U134 ( .A1(D[26]), .A2(n1420), .B1(C[26]), .B2(n1414), .ZN(n192) );
  NAND4_X1 U135 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U136 ( .A1(B[46]), .A2(n1410), .B1(A[46]), .B2(n1404), .ZN(n103) );
  AOI22_X1 U137 ( .A1(D[46]), .A2(n1422), .B1(C[46]), .B2(n1416), .ZN(n104) );
  AOI22_X1 U138 ( .A1(H[46]), .A2(n1446), .B1(G[46]), .B2(n1440), .ZN(n106) );
  NAND4_X1 U139 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U140 ( .A1(B[41]), .A2(n1409), .B1(A[41]), .B2(n1403), .ZN(n123) );
  AOI22_X1 U141 ( .A1(D[41]), .A2(n1421), .B1(C[41]), .B2(n1415), .ZN(n124) );
  AOI22_X1 U142 ( .A1(H[41]), .A2(n1445), .B1(G[41]), .B2(n1439), .ZN(n126) );
  NAND4_X1 U143 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U144 ( .A1(B[34]), .A2(n1409), .B1(A[34]), .B2(n1403), .ZN(n155) );
  AOI22_X1 U145 ( .A1(D[34]), .A2(n1421), .B1(C[34]), .B2(n1415), .ZN(n156) );
  AOI22_X1 U146 ( .A1(H[34]), .A2(n1445), .B1(G[34]), .B2(n1439), .ZN(n158) );
  NAND4_X1 U147 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U148 ( .A1(B[37]), .A2(n1409), .B1(A[37]), .B2(n1403), .ZN(n143) );
  AOI22_X1 U149 ( .A1(D[37]), .A2(n1421), .B1(C[37]), .B2(n1415), .ZN(n144) );
  AOI22_X1 U150 ( .A1(H[37]), .A2(n1445), .B1(G[37]), .B2(n1439), .ZN(n146) );
  NAND4_X1 U151 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U152 ( .A1(H[26]), .A2(n1444), .B1(G[26]), .B2(n1438), .ZN(n194) );
  AOI22_X1 U153 ( .A1(B[26]), .A2(n1408), .B1(A[26]), .B2(n1402), .ZN(n191) );
  AOI22_X1 U154 ( .A1(F[26]), .A2(n1432), .B1(E[26]), .B2(n1426), .ZN(n193) );
  NAND4_X1 U155 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U156 ( .A1(H[23]), .A2(n1444), .B1(G[23]), .B2(n1438), .ZN(n206) );
  AOI22_X1 U157 ( .A1(B[23]), .A2(n1408), .B1(A[23]), .B2(n1402), .ZN(n203) );
  AOI22_X1 U158 ( .A1(D[23]), .A2(n1420), .B1(C[23]), .B2(n1414), .ZN(n204) );
  NAND4_X1 U159 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U160 ( .A1(B[24]), .A2(n1408), .B1(A[24]), .B2(n1402), .ZN(n199) );
  AOI22_X1 U161 ( .A1(H[24]), .A2(n1444), .B1(G[24]), .B2(n1438), .ZN(n202) );
  AOI22_X1 U162 ( .A1(F[24]), .A2(n1432), .B1(E[24]), .B2(n1426), .ZN(n201) );
  NAND4_X1 U163 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U164 ( .A1(B[25]), .A2(n1408), .B1(A[25]), .B2(n1402), .ZN(n195) );
  AOI22_X1 U165 ( .A1(H[25]), .A2(n1444), .B1(G[25]), .B2(n1438), .ZN(n198) );
  AOI22_X1 U166 ( .A1(F[25]), .A2(n1432), .B1(E[25]), .B2(n1426), .ZN(n197) );
  NAND4_X1 U167 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U168 ( .A1(B[29]), .A2(n1408), .B1(A[29]), .B2(n1402), .ZN(n179) );
  AOI22_X1 U169 ( .A1(H[29]), .A2(n1444), .B1(G[29]), .B2(n1438), .ZN(n182) );
  AOI22_X1 U170 ( .A1(D[29]), .A2(n1420), .B1(C[29]), .B2(n1414), .ZN(n180) );
  NAND4_X1 U171 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U172 ( .A1(B[32]), .A2(n1409), .B1(A[32]), .B2(n1403), .ZN(n163) );
  AOI22_X1 U173 ( .A1(D[32]), .A2(n1421), .B1(C[32]), .B2(n1415), .ZN(n164) );
  AOI22_X1 U174 ( .A1(H[32]), .A2(n1445), .B1(G[32]), .B2(n1439), .ZN(n166) );
  NAND4_X1 U175 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U176 ( .A1(B[36]), .A2(n1409), .B1(A[36]), .B2(n1403), .ZN(n147) );
  AOI22_X1 U177 ( .A1(D[36]), .A2(n1421), .B1(C[36]), .B2(n1415), .ZN(n148) );
  AOI22_X1 U178 ( .A1(H[36]), .A2(n1445), .B1(G[36]), .B2(n1439), .ZN(n150) );
  NAND4_X1 U179 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U180 ( .A1(B[39]), .A2(n1409), .B1(A[39]), .B2(n1403), .ZN(n135) );
  AOI22_X1 U181 ( .A1(D[39]), .A2(n1421), .B1(C[39]), .B2(n1415), .ZN(n136) );
  AOI22_X1 U182 ( .A1(H[39]), .A2(n1445), .B1(G[39]), .B2(n1439), .ZN(n138) );
  NAND4_X1 U183 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U184 ( .A1(B[40]), .A2(n1409), .B1(A[40]), .B2(n1403), .ZN(n127) );
  AOI22_X1 U185 ( .A1(D[40]), .A2(n1421), .B1(C[40]), .B2(n1415), .ZN(n128) );
  AOI22_X1 U186 ( .A1(H[40]), .A2(n1445), .B1(G[40]), .B2(n1439), .ZN(n130) );
  NAND4_X1 U187 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U188 ( .A1(D[22]), .A2(n1420), .B1(C[22]), .B2(n1414), .ZN(n208) );
  AOI22_X1 U189 ( .A1(H[22]), .A2(n1444), .B1(G[22]), .B2(n1438), .ZN(n210) );
  AOI22_X1 U190 ( .A1(B[22]), .A2(n1408), .B1(A[22]), .B2(n1402), .ZN(n207) );
  NAND4_X1 U191 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U192 ( .A1(B[55]), .A2(n1411), .B1(A[55]), .B2(n1405), .ZN(n63) );
  AOI22_X1 U193 ( .A1(D[55]), .A2(n1423), .B1(C[55]), .B2(n1417), .ZN(n64) );
  AOI22_X1 U194 ( .A1(H[55]), .A2(n1447), .B1(G[55]), .B2(n1441), .ZN(n66) );
  NAND4_X1 U195 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U196 ( .A1(B[62]), .A2(n1411), .B1(A[62]), .B2(n1405), .ZN(n31) );
  AOI22_X1 U197 ( .A1(D[62]), .A2(n1423), .B1(C[62]), .B2(n1417), .ZN(n32) );
  AOI22_X1 U198 ( .A1(H[62]), .A2(n1447), .B1(G[62]), .B2(n1441), .ZN(n34) );
  NAND4_X1 U199 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U200 ( .A1(B[31]), .A2(n1409), .B1(A[31]), .B2(n1403), .ZN(n167) );
  AOI22_X1 U201 ( .A1(D[31]), .A2(n1421), .B1(C[31]), .B2(n1415), .ZN(n168) );
  AOI22_X1 U202 ( .A1(H[31]), .A2(n1445), .B1(G[31]), .B2(n1439), .ZN(n170) );
  NAND4_X1 U203 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U204 ( .A1(H[28]), .A2(n1444), .B1(G[28]), .B2(n1438), .ZN(n186) );
  AOI22_X1 U205 ( .A1(B[28]), .A2(n1408), .B1(A[28]), .B2(n1402), .ZN(n183) );
  AOI22_X1 U206 ( .A1(F[28]), .A2(n1432), .B1(E[28]), .B2(n1426), .ZN(n185) );
  NAND4_X1 U207 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U208 ( .A1(B[38]), .A2(n1409), .B1(A[38]), .B2(n1403), .ZN(n139) );
  AOI22_X1 U209 ( .A1(D[38]), .A2(n1421), .B1(C[38]), .B2(n1415), .ZN(n140) );
  AOI22_X1 U210 ( .A1(H[38]), .A2(n1445), .B1(G[38]), .B2(n1439), .ZN(n142) );
  NAND4_X1 U211 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U212 ( .A1(B[33]), .A2(n1409), .B1(A[33]), .B2(n1403), .ZN(n159) );
  AOI22_X1 U213 ( .A1(D[33]), .A2(n1421), .B1(C[33]), .B2(n1415), .ZN(n160) );
  AOI22_X1 U214 ( .A1(H[33]), .A2(n1445), .B1(G[33]), .B2(n1439), .ZN(n162) );
  AOI22_X1 U215 ( .A1(F[60]), .A2(n1435), .B1(E[60]), .B2(n1429), .ZN(n41) );
  AOI22_X1 U216 ( .A1(F[56]), .A2(n1435), .B1(E[56]), .B2(n1429), .ZN(n61) );
  AOI22_X1 U217 ( .A1(F[52]), .A2(n1434), .B1(E[52]), .B2(n1428), .ZN(n77) );
  AOI22_X1 U218 ( .A1(F[48]), .A2(n1434), .B1(E[48]), .B2(n1428), .ZN(n97) );
  NAND4_X1 U219 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U220 ( .A1(B[57]), .A2(n1411), .B1(A[57]), .B2(n1405), .ZN(n55) );
  AOI22_X1 U221 ( .A1(D[57]), .A2(n1423), .B1(C[57]), .B2(n1417), .ZN(n56) );
  AOI22_X1 U222 ( .A1(H[57]), .A2(n1447), .B1(G[57]), .B2(n1441), .ZN(n58) );
  NAND4_X1 U223 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U224 ( .A1(B[27]), .A2(n1408), .B1(A[27]), .B2(n1402), .ZN(n187) );
  AOI22_X1 U225 ( .A1(H[27]), .A2(n1444), .B1(G[27]), .B2(n1438), .ZN(n190) );
  AOI22_X1 U226 ( .A1(F[27]), .A2(n1432), .B1(E[27]), .B2(n1426), .ZN(n189) );
  NAND4_X1 U227 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U228 ( .A1(B[44]), .A2(n1410), .B1(A[44]), .B2(n1404), .ZN(n111) );
  AOI22_X1 U229 ( .A1(D[44]), .A2(n1422), .B1(C[44]), .B2(n1416), .ZN(n112) );
  AOI22_X1 U230 ( .A1(H[44]), .A2(n1446), .B1(G[44]), .B2(n1440), .ZN(n114) );
  NAND4_X1 U231 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U232 ( .A1(B[56]), .A2(n1411), .B1(A[56]), .B2(n1405), .ZN(n59) );
  AOI22_X1 U233 ( .A1(D[56]), .A2(n1423), .B1(C[56]), .B2(n1417), .ZN(n60) );
  AOI22_X1 U234 ( .A1(H[56]), .A2(n1447), .B1(G[56]), .B2(n1441), .ZN(n62) );
  NAND4_X1 U235 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U236 ( .A1(B[58]), .A2(n1411), .B1(A[58]), .B2(n1405), .ZN(n51) );
  AOI22_X1 U237 ( .A1(D[58]), .A2(n1423), .B1(C[58]), .B2(n1417), .ZN(n52) );
  AOI22_X1 U238 ( .A1(H[58]), .A2(n1447), .B1(G[58]), .B2(n1441), .ZN(n54) );
  NAND4_X1 U239 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U240 ( .A1(B[54]), .A2(n1411), .B1(A[54]), .B2(n1405), .ZN(n67) );
  AOI22_X1 U241 ( .A1(D[54]), .A2(n1423), .B1(C[54]), .B2(n1417), .ZN(n68) );
  AOI22_X1 U242 ( .A1(H[54]), .A2(n1447), .B1(G[54]), .B2(n1441), .ZN(n70) );
  NAND4_X1 U243 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U244 ( .A1(B[59]), .A2(n1411), .B1(A[59]), .B2(n1405), .ZN(n47) );
  AOI22_X1 U245 ( .A1(D[59]), .A2(n1423), .B1(C[59]), .B2(n1417), .ZN(n48) );
  AOI22_X1 U246 ( .A1(H[59]), .A2(n1447), .B1(G[59]), .B2(n1441), .ZN(n50) );
  NAND4_X1 U247 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U248 ( .A1(B[60]), .A2(n1411), .B1(A[60]), .B2(n1405), .ZN(n39) );
  AOI22_X1 U249 ( .A1(D[60]), .A2(n1423), .B1(C[60]), .B2(n1417), .ZN(n40) );
  AOI22_X1 U250 ( .A1(H[60]), .A2(n1447), .B1(G[60]), .B2(n1441), .ZN(n42) );
  NAND4_X1 U251 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U252 ( .A1(B[63]), .A2(n1411), .B1(A[63]), .B2(n1405), .ZN(n27) );
  AOI22_X1 U253 ( .A1(D[63]), .A2(n1423), .B1(C[63]), .B2(n1417), .ZN(n28) );
  AOI22_X1 U254 ( .A1(H[63]), .A2(n1447), .B1(G[63]), .B2(n1441), .ZN(n30) );
  AOI22_X1 U255 ( .A1(F[46]), .A2(n1434), .B1(E[46]), .B2(n1428), .ZN(n105) );
  AOI22_X1 U256 ( .A1(F[34]), .A2(n1433), .B1(E[34]), .B2(n1427), .ZN(n157) );
  NAND4_X1 U257 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U258 ( .A1(B[61]), .A2(n1411), .B1(A[61]), .B2(n1405), .ZN(n35) );
  AOI22_X1 U259 ( .A1(D[61]), .A2(n1423), .B1(C[61]), .B2(n1417), .ZN(n36) );
  AOI22_X1 U260 ( .A1(H[61]), .A2(n1447), .B1(G[61]), .B2(n1441), .ZN(n38) );
  NAND4_X1 U261 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U262 ( .A1(B[0]), .A2(n1407), .B1(A[0]), .B2(n1401), .ZN(n263) );
  AOI22_X1 U263 ( .A1(D[0]), .A2(n1419), .B1(C[0]), .B2(n1413), .ZN(n264) );
  AOI22_X1 U264 ( .A1(F[0]), .A2(n1431), .B1(E[0]), .B2(n1425), .ZN(n265) );
  AOI22_X1 U265 ( .A1(H[5]), .A2(n1447), .B1(G[5]), .B2(n1441), .ZN(n46) );
  AOI22_X1 U266 ( .A1(H[13]), .A2(n1443), .B1(G[13]), .B2(n1437), .ZN(n250) );
  AOI22_X1 U267 ( .A1(H[17]), .A2(n1443), .B1(G[17]), .B2(n1437), .ZN(n234) );
  AOI22_X1 U268 ( .A1(H[21]), .A2(n1444), .B1(G[21]), .B2(n1438), .ZN(n214) );
  AOI22_X1 U269 ( .A1(H[9]), .A2(n1448), .B1(G[9]), .B2(n1442), .ZN(n6) );
  AOI22_X1 U270 ( .A1(H[7]), .A2(n1448), .B1(G[7]), .B2(n1442), .ZN(n22) );
  AOI22_X1 U271 ( .A1(H[11]), .A2(n1443), .B1(G[11]), .B2(n1437), .ZN(n258) );
  AOI22_X1 U272 ( .A1(H[15]), .A2(n1443), .B1(G[15]), .B2(n1437), .ZN(n242) );
  AOI22_X1 U273 ( .A1(H[19]), .A2(n1443), .B1(G[19]), .B2(n1437), .ZN(n226) );
  AOI22_X1 U274 ( .A1(H[3]), .A2(n1445), .B1(G[3]), .B2(n1439), .ZN(n134) );
  AOI22_X1 U275 ( .A1(H[4]), .A2(n1446), .B1(G[4]), .B2(n1440), .ZN(n90) );
  AOI22_X1 U276 ( .A1(H[16]), .A2(n1443), .B1(G[16]), .B2(n1437), .ZN(n238) );
  AOI22_X1 U277 ( .A1(H[20]), .A2(n1444), .B1(G[20]), .B2(n1438), .ZN(n218) );
  AOI22_X1 U278 ( .A1(H[12]), .A2(n1443), .B1(G[12]), .B2(n1437), .ZN(n254) );
  AOI22_X1 U279 ( .A1(H[8]), .A2(n1448), .B1(G[8]), .B2(n1442), .ZN(n18) );
  AOI22_X1 U280 ( .A1(H[6]), .A2(n1448), .B1(G[6]), .B2(n1442), .ZN(n26) );
  AOI22_X1 U281 ( .A1(H[10]), .A2(n1443), .B1(G[10]), .B2(n1437), .ZN(n262) );
  AOI22_X1 U282 ( .A1(H[14]), .A2(n1443), .B1(G[14]), .B2(n1437), .ZN(n246) );
  AOI22_X1 U283 ( .A1(H[18]), .A2(n1443), .B1(G[18]), .B2(n1437), .ZN(n230) );
  AOI22_X1 U284 ( .A1(H[2]), .A2(n1444), .B1(G[2]), .B2(n1438), .ZN(n178) );
  AOI22_X1 U285 ( .A1(H[1]), .A2(n1443), .B1(G[1]), .B2(n1437), .ZN(n222) );
  NAND4_X1 U286 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U287 ( .A1(B[4]), .A2(n1410), .B1(A[4]), .B2(n1404), .ZN(n87) );
  AOI22_X1 U288 ( .A1(D[4]), .A2(n1422), .B1(C[4]), .B2(n1416), .ZN(n88) );
  AOI22_X1 U289 ( .A1(F[4]), .A2(n1434), .B1(E[4]), .B2(n1428), .ZN(n89) );
  NAND4_X1 U290 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U291 ( .A1(B[5]), .A2(n1411), .B1(A[5]), .B2(n1405), .ZN(n43) );
  AOI22_X1 U292 ( .A1(D[5]), .A2(n1423), .B1(C[5]), .B2(n1417), .ZN(n44) );
  AOI22_X1 U293 ( .A1(F[5]), .A2(n1435), .B1(E[5]), .B2(n1429), .ZN(n45) );
  NAND4_X1 U294 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U295 ( .A1(B[13]), .A2(n1407), .B1(A[13]), .B2(n1401), .ZN(n247) );
  AOI22_X1 U296 ( .A1(D[13]), .A2(n1419), .B1(C[13]), .B2(n1413), .ZN(n248) );
  AOI22_X1 U297 ( .A1(F[13]), .A2(n1431), .B1(E[13]), .B2(n1425), .ZN(n249) );
  NAND4_X1 U298 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U299 ( .A1(B[17]), .A2(n1407), .B1(A[17]), .B2(n1401), .ZN(n231) );
  AOI22_X1 U300 ( .A1(D[17]), .A2(n1419), .B1(C[17]), .B2(n1413), .ZN(n232) );
  AOI22_X1 U301 ( .A1(F[17]), .A2(n1431), .B1(E[17]), .B2(n1425), .ZN(n233) );
  NAND4_X1 U302 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U303 ( .A1(B[16]), .A2(n1407), .B1(A[16]), .B2(n1401), .ZN(n235) );
  AOI22_X1 U304 ( .A1(D[16]), .A2(n1419), .B1(C[16]), .B2(n1413), .ZN(n236) );
  AOI22_X1 U305 ( .A1(F[16]), .A2(n1431), .B1(E[16]), .B2(n1425), .ZN(n237) );
  NAND4_X1 U306 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U307 ( .A1(B[12]), .A2(n1407), .B1(A[12]), .B2(n1401), .ZN(n251) );
  AOI22_X1 U308 ( .A1(D[12]), .A2(n1419), .B1(C[12]), .B2(n1413), .ZN(n252) );
  AOI22_X1 U309 ( .A1(F[12]), .A2(n1431), .B1(E[12]), .B2(n1425), .ZN(n253) );
  NAND4_X1 U310 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U311 ( .A1(B[21]), .A2(n1408), .B1(A[21]), .B2(n1402), .ZN(n211) );
  AOI22_X1 U312 ( .A1(D[21]), .A2(n1420), .B1(C[21]), .B2(n1414), .ZN(n212) );
  AOI22_X1 U313 ( .A1(F[21]), .A2(n1432), .B1(E[21]), .B2(n1426), .ZN(n213) );
  NAND4_X1 U314 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U315 ( .A1(B[8]), .A2(n1412), .B1(A[8]), .B2(n1406), .ZN(n15) );
  AOI22_X1 U316 ( .A1(D[8]), .A2(n1424), .B1(C[8]), .B2(n1418), .ZN(n16) );
  AOI22_X1 U317 ( .A1(F[8]), .A2(n1436), .B1(E[8]), .B2(n1430), .ZN(n17) );
  NAND4_X1 U318 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U319 ( .A1(B[9]), .A2(n1412), .B1(A[9]), .B2(n1406), .ZN(n3) );
  AOI22_X1 U320 ( .A1(D[9]), .A2(n1424), .B1(C[9]), .B2(n1418), .ZN(n4) );
  AOI22_X1 U321 ( .A1(F[9]), .A2(n1436), .B1(E[9]), .B2(n1430), .ZN(n5) );
  NAND4_X1 U322 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U323 ( .A1(B[7]), .A2(n1412), .B1(A[7]), .B2(n1406), .ZN(n19) );
  AOI22_X1 U324 ( .A1(D[7]), .A2(n1424), .B1(C[7]), .B2(n1418), .ZN(n20) );
  AOI22_X1 U325 ( .A1(F[7]), .A2(n1436), .B1(E[7]), .B2(n1430), .ZN(n21) );
  NAND4_X1 U326 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U327 ( .A1(B[11]), .A2(n1407), .B1(A[11]), .B2(n1401), .ZN(n255) );
  AOI22_X1 U328 ( .A1(D[11]), .A2(n1419), .B1(C[11]), .B2(n1413), .ZN(n256) );
  AOI22_X1 U329 ( .A1(F[11]), .A2(n1431), .B1(E[11]), .B2(n1425), .ZN(n257) );
  NAND4_X1 U330 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U331 ( .A1(B[15]), .A2(n1407), .B1(A[15]), .B2(n1401), .ZN(n239) );
  AOI22_X1 U332 ( .A1(D[15]), .A2(n1419), .B1(C[15]), .B2(n1413), .ZN(n240) );
  AOI22_X1 U333 ( .A1(F[15]), .A2(n1431), .B1(E[15]), .B2(n1425), .ZN(n241) );
  NAND4_X1 U334 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U335 ( .A1(B[3]), .A2(n1409), .B1(A[3]), .B2(n1403), .ZN(n131) );
  AOI22_X1 U336 ( .A1(D[3]), .A2(n1421), .B1(C[3]), .B2(n1415), .ZN(n132) );
  AOI22_X1 U337 ( .A1(F[3]), .A2(n1433), .B1(E[3]), .B2(n1427), .ZN(n133) );
  NAND4_X1 U338 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U339 ( .A1(B[20]), .A2(n1408), .B1(A[20]), .B2(n1402), .ZN(n215) );
  AOI22_X1 U340 ( .A1(D[20]), .A2(n1420), .B1(C[20]), .B2(n1414), .ZN(n216) );
  AOI22_X1 U341 ( .A1(F[20]), .A2(n1432), .B1(E[20]), .B2(n1426), .ZN(n217) );
  NAND4_X1 U342 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U343 ( .A1(B[19]), .A2(n1407), .B1(A[19]), .B2(n1401), .ZN(n223) );
  AOI22_X1 U344 ( .A1(D[19]), .A2(n1419), .B1(C[19]), .B2(n1413), .ZN(n224) );
  AOI22_X1 U345 ( .A1(F[19]), .A2(n1431), .B1(E[19]), .B2(n1425), .ZN(n225) );
  NAND4_X1 U346 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U347 ( .A1(B[6]), .A2(n1412), .B1(A[6]), .B2(n1406), .ZN(n23) );
  AOI22_X1 U348 ( .A1(D[6]), .A2(n1424), .B1(C[6]), .B2(n1418), .ZN(n24) );
  AOI22_X1 U349 ( .A1(F[6]), .A2(n1436), .B1(E[6]), .B2(n1430), .ZN(n25) );
  NAND4_X1 U350 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U351 ( .A1(B[10]), .A2(n1407), .B1(A[10]), .B2(n1401), .ZN(n259) );
  AOI22_X1 U352 ( .A1(D[10]), .A2(n1419), .B1(C[10]), .B2(n1413), .ZN(n260) );
  AOI22_X1 U353 ( .A1(F[10]), .A2(n1431), .B1(E[10]), .B2(n1425), .ZN(n261) );
  NAND4_X1 U354 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U355 ( .A1(B[14]), .A2(n1407), .B1(A[14]), .B2(n1401), .ZN(n243) );
  AOI22_X1 U356 ( .A1(D[14]), .A2(n1419), .B1(C[14]), .B2(n1413), .ZN(n244) );
  AOI22_X1 U357 ( .A1(F[14]), .A2(n1431), .B1(E[14]), .B2(n1425), .ZN(n245) );
  NAND4_X1 U358 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U359 ( .A1(B[18]), .A2(n1407), .B1(A[18]), .B2(n1401), .ZN(n227) );
  AOI22_X1 U360 ( .A1(D[18]), .A2(n1419), .B1(C[18]), .B2(n1413), .ZN(n228) );
  AOI22_X1 U361 ( .A1(F[18]), .A2(n1431), .B1(E[18]), .B2(n1425), .ZN(n229) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1408), .B1(A[2]), .B2(n1402), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1420), .B1(C[2]), .B2(n1414), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1432), .B1(E[2]), .B2(n1426), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1407), .B1(A[1]), .B2(n1401), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1419), .B1(C[1]), .B2(n1413), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1431), .B1(E[1]), .B2(n1425), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1443), .B1(G[0]), .B2(n1437), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1406) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1412) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1418) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1424) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1430) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1436) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1442) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1448) );
endmodule


module MUX81_GENERIC_NBIT64_4 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446;

  BUF_X1 U1 ( .A(n13), .Z(n1404) );
  BUF_X1 U2 ( .A(n12), .Z(n1410) );
  BUF_X1 U3 ( .A(n8), .Z(n1434) );
  BUF_X1 U4 ( .A(n10), .Z(n1422) );
  BUF_X1 U5 ( .A(n13), .Z(n1406) );
  BUF_X1 U6 ( .A(n13), .Z(n1405) );
  BUF_X1 U7 ( .A(n13), .Z(n1407) );
  BUF_X1 U8 ( .A(n12), .Z(n1412) );
  BUF_X1 U9 ( .A(n12), .Z(n1411) );
  BUF_X1 U10 ( .A(n12), .Z(n1413) );
  BUF_X1 U11 ( .A(n8), .Z(n1435) );
  BUF_X1 U12 ( .A(n10), .Z(n1424) );
  BUF_X1 U13 ( .A(n8), .Z(n1436) );
  BUF_X1 U14 ( .A(n10), .Z(n1425) );
  BUF_X1 U15 ( .A(n10), .Z(n1423) );
  BUF_X1 U16 ( .A(n8), .Z(n1437) );
  BUF_X1 U17 ( .A(n11), .Z(n1418) );
  BUF_X1 U18 ( .A(n11), .Z(n1416) );
  BUF_X1 U19 ( .A(n11), .Z(n1417) );
  BUF_X1 U20 ( .A(n11), .Z(n1415) );
  BUF_X1 U21 ( .A(n13), .Z(n1403) );
  BUF_X1 U22 ( .A(n11), .Z(n1419) );
  BUF_X1 U23 ( .A(n7), .Z(n1439) );
  BUF_X1 U24 ( .A(n7), .Z(n1441) );
  BUF_X1 U25 ( .A(n9), .Z(n1430) );
  BUF_X1 U26 ( .A(n7), .Z(n1442) );
  BUF_X1 U27 ( .A(n7), .Z(n1440) );
  BUF_X1 U28 ( .A(n9), .Z(n1431) );
  BUF_X1 U29 ( .A(n9), .Z(n1428) );
  BUF_X1 U30 ( .A(n9), .Z(n1429) );
  BUF_X1 U31 ( .A(n9), .Z(n1427) );
  BUF_X1 U32 ( .A(n7), .Z(n1443) );
  BUF_X1 U33 ( .A(n14), .Z(n1400) );
  BUF_X1 U34 ( .A(n14), .Z(n1398) );
  BUF_X1 U35 ( .A(n14), .Z(n1399) );
  BUF_X1 U36 ( .A(n12), .Z(n1409) );
  BUF_X1 U37 ( .A(n14), .Z(n1397) );
  BUF_X1 U38 ( .A(n14), .Z(n1401) );
  BUF_X1 U39 ( .A(n8), .Z(n1433) );
  BUF_X1 U40 ( .A(n10), .Z(n1421) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1445), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1446), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1446), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1446), .A2(n1445), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1445) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1446) );
  NOR3_X1 U47 ( .A1(n1446), .A2(SEL[2]), .A3(n1445), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1445), .A3(SEL[2]), .ZN(n9) );
  AOI22_X1 U51 ( .A1(F[43]), .A2(n1430), .B1(E[43]), .B2(n1424), .ZN(n117) );
  AOI22_X1 U52 ( .A1(F[62]), .A2(n1431), .B1(E[62]), .B2(n1425), .ZN(n33) );
  AOI22_X1 U53 ( .A1(F[57]), .A2(n1431), .B1(E[57]), .B2(n1425), .ZN(n57) );
  AOI22_X1 U54 ( .A1(F[53]), .A2(n1431), .B1(E[53]), .B2(n1425), .ZN(n73) );
  AOI22_X1 U55 ( .A1(F[61]), .A2(n1431), .B1(E[61]), .B2(n1425), .ZN(n37) );
  NAND4_X1 U56 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U57 ( .A1(H[25]), .A2(n1440), .B1(G[25]), .B2(n1434), .ZN(n198) );
  AOI22_X1 U58 ( .A1(B[25]), .A2(n1404), .B1(A[25]), .B2(n1398), .ZN(n195) );
  AOI22_X1 U59 ( .A1(F[25]), .A2(n1428), .B1(E[25]), .B2(n1422), .ZN(n197) );
  NAND4_X1 U60 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U61 ( .A1(B[41]), .A2(n1405), .B1(A[41]), .B2(n1399), .ZN(n123) );
  AOI22_X1 U62 ( .A1(D[41]), .A2(n1417), .B1(C[41]), .B2(n1411), .ZN(n124) );
  AOI22_X1 U63 ( .A1(H[41]), .A2(n1441), .B1(G[41]), .B2(n1435), .ZN(n126) );
  NAND4_X1 U64 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U65 ( .A1(B[47]), .A2(n1406), .B1(A[47]), .B2(n1400), .ZN(n99) );
  AOI22_X1 U66 ( .A1(D[47]), .A2(n1418), .B1(C[47]), .B2(n1412), .ZN(n100) );
  AOI22_X1 U67 ( .A1(H[47]), .A2(n1442), .B1(G[47]), .B2(n1436), .ZN(n102) );
  NAND4_X1 U68 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U69 ( .A1(B[39]), .A2(n1405), .B1(A[39]), .B2(n1399), .ZN(n135) );
  AOI22_X1 U70 ( .A1(D[39]), .A2(n1417), .B1(C[39]), .B2(n1411), .ZN(n136) );
  AOI22_X1 U71 ( .A1(H[39]), .A2(n1441), .B1(G[39]), .B2(n1435), .ZN(n138) );
  NAND4_X1 U72 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U73 ( .A1(B[46]), .A2(n1406), .B1(A[46]), .B2(n1400), .ZN(n103) );
  AOI22_X1 U74 ( .A1(D[46]), .A2(n1418), .B1(C[46]), .B2(n1412), .ZN(n104) );
  AOI22_X1 U75 ( .A1(H[46]), .A2(n1442), .B1(G[46]), .B2(n1436), .ZN(n106) );
  NAND4_X1 U76 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U77 ( .A1(B[54]), .A2(n1407), .B1(A[54]), .B2(n1401), .ZN(n67) );
  AOI22_X1 U78 ( .A1(D[54]), .A2(n1419), .B1(C[54]), .B2(n1413), .ZN(n68) );
  AOI22_X1 U79 ( .A1(H[54]), .A2(n1443), .B1(G[54]), .B2(n1437), .ZN(n70) );
  NAND4_X1 U80 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U81 ( .A1(B[57]), .A2(n1407), .B1(A[57]), .B2(n1401), .ZN(n55) );
  AOI22_X1 U82 ( .A1(D[57]), .A2(n1419), .B1(C[57]), .B2(n1413), .ZN(n56) );
  AOI22_X1 U83 ( .A1(H[57]), .A2(n1443), .B1(G[57]), .B2(n1437), .ZN(n58) );
  NAND4_X1 U84 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U85 ( .A1(B[42]), .A2(n1406), .B1(A[42]), .B2(n1400), .ZN(n119) );
  AOI22_X1 U86 ( .A1(D[42]), .A2(n1418), .B1(C[42]), .B2(n1412), .ZN(n120) );
  AOI22_X1 U87 ( .A1(H[42]), .A2(n1442), .B1(G[42]), .B2(n1436), .ZN(n122) );
  AOI22_X1 U88 ( .A1(F[29]), .A2(n1428), .B1(E[29]), .B2(n1422), .ZN(n181) );
  AOI22_X1 U89 ( .A1(F[28]), .A2(n1428), .B1(E[28]), .B2(n1422), .ZN(n185) );
  AOI22_X1 U90 ( .A1(F[31]), .A2(n1429), .B1(E[31]), .B2(n1423), .ZN(n169) );
  AOI22_X1 U91 ( .A1(F[35]), .A2(n1429), .B1(E[35]), .B2(n1423), .ZN(n153) );
  AOI22_X1 U92 ( .A1(F[32]), .A2(n1429), .B1(E[32]), .B2(n1423), .ZN(n165) );
  AOI22_X1 U93 ( .A1(F[33]), .A2(n1429), .B1(E[33]), .B2(n1423), .ZN(n161) );
  AOI22_X1 U94 ( .A1(F[30]), .A2(n1428), .B1(E[30]), .B2(n1422), .ZN(n173) );
  AOI22_X1 U95 ( .A1(F[39]), .A2(n1429), .B1(E[39]), .B2(n1423), .ZN(n137) );
  AOI22_X1 U96 ( .A1(F[37]), .A2(n1429), .B1(E[37]), .B2(n1423), .ZN(n145) );
  AOI22_X1 U97 ( .A1(F[40]), .A2(n1429), .B1(E[40]), .B2(n1423), .ZN(n129) );
  AOI22_X1 U98 ( .A1(F[24]), .A2(n1428), .B1(E[24]), .B2(n1422), .ZN(n201) );
  AOI22_X1 U99 ( .A1(F[41]), .A2(n1429), .B1(E[41]), .B2(n1423), .ZN(n125) );
  AOI22_X1 U100 ( .A1(F[45]), .A2(n1430), .B1(E[45]), .B2(n1424), .ZN(n109) );
  AOI22_X1 U101 ( .A1(F[44]), .A2(n1430), .B1(E[44]), .B2(n1424), .ZN(n113) );
  AOI22_X1 U102 ( .A1(F[34]), .A2(n1429), .B1(E[34]), .B2(n1423), .ZN(n157) );
  AOI22_X1 U103 ( .A1(F[47]), .A2(n1430), .B1(E[47]), .B2(n1424), .ZN(n101) );
  AOI22_X1 U104 ( .A1(F[51]), .A2(n1430), .B1(E[51]), .B2(n1424), .ZN(n81) );
  AOI22_X1 U105 ( .A1(F[49]), .A2(n1430), .B1(E[49]), .B2(n1424), .ZN(n93) );
  AOI22_X1 U106 ( .A1(F[52]), .A2(n1430), .B1(E[52]), .B2(n1424), .ZN(n77) );
  AOI22_X1 U107 ( .A1(F[26]), .A2(n1428), .B1(E[26]), .B2(n1422), .ZN(n193) );
  AOI22_X1 U108 ( .A1(F[55]), .A2(n1431), .B1(E[55]), .B2(n1425), .ZN(n65) );
  AOI22_X1 U109 ( .A1(F[27]), .A2(n1428), .B1(E[27]), .B2(n1422), .ZN(n189) );
  AOI22_X1 U110 ( .A1(F[58]), .A2(n1431), .B1(E[58]), .B2(n1425), .ZN(n53) );
  AOI22_X1 U111 ( .A1(F[59]), .A2(n1431), .B1(E[59]), .B2(n1425), .ZN(n49) );
  AOI22_X1 U112 ( .A1(F[60]), .A2(n1431), .B1(E[60]), .B2(n1425), .ZN(n41) );
  AOI22_X1 U113 ( .A1(F[63]), .A2(n1431), .B1(E[63]), .B2(n1425), .ZN(n29) );
  NAND4_X1 U114 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U115 ( .A1(B[35]), .A2(n1405), .B1(A[35]), .B2(n1399), .ZN(n151) );
  AOI22_X1 U116 ( .A1(D[35]), .A2(n1417), .B1(C[35]), .B2(n1411), .ZN(n152) );
  AOI22_X1 U117 ( .A1(H[35]), .A2(n1441), .B1(G[35]), .B2(n1435), .ZN(n154) );
  AOI22_X1 U118 ( .A1(D[25]), .A2(n1416), .B1(C[25]), .B2(n1410), .ZN(n196) );
  NAND4_X1 U119 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U120 ( .A1(B[58]), .A2(n1407), .B1(A[58]), .B2(n1401), .ZN(n51) );
  AOI22_X1 U121 ( .A1(D[58]), .A2(n1419), .B1(C[58]), .B2(n1413), .ZN(n52) );
  AOI22_X1 U122 ( .A1(H[58]), .A2(n1443), .B1(G[58]), .B2(n1437), .ZN(n54) );
  NAND4_X1 U123 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U124 ( .A1(B[53]), .A2(n1407), .B1(A[53]), .B2(n1401), .ZN(n71) );
  AOI22_X1 U125 ( .A1(D[53]), .A2(n1419), .B1(C[53]), .B2(n1413), .ZN(n72) );
  AOI22_X1 U126 ( .A1(H[53]), .A2(n1443), .B1(G[53]), .B2(n1437), .ZN(n74) );
  NAND4_X1 U127 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U128 ( .A1(B[44]), .A2(n1406), .B1(A[44]), .B2(n1400), .ZN(n111) );
  AOI22_X1 U129 ( .A1(D[44]), .A2(n1418), .B1(C[44]), .B2(n1412), .ZN(n112) );
  AOI22_X1 U130 ( .A1(H[44]), .A2(n1442), .B1(G[44]), .B2(n1436), .ZN(n114) );
  NAND4_X1 U131 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U132 ( .A1(B[45]), .A2(n1406), .B1(A[45]), .B2(n1400), .ZN(n107) );
  AOI22_X1 U133 ( .A1(D[45]), .A2(n1418), .B1(C[45]), .B2(n1412), .ZN(n108) );
  AOI22_X1 U134 ( .A1(H[45]), .A2(n1442), .B1(G[45]), .B2(n1436), .ZN(n110) );
  NAND4_X1 U135 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U136 ( .A1(B[49]), .A2(n1406), .B1(A[49]), .B2(n1400), .ZN(n91) );
  AOI22_X1 U137 ( .A1(D[49]), .A2(n1418), .B1(C[49]), .B2(n1412), .ZN(n92) );
  AOI22_X1 U138 ( .A1(H[49]), .A2(n1442), .B1(G[49]), .B2(n1436), .ZN(n94) );
  NAND4_X1 U139 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U140 ( .A1(H[27]), .A2(n1440), .B1(G[27]), .B2(n1434), .ZN(n190) );
  AOI22_X1 U141 ( .A1(B[27]), .A2(n1404), .B1(A[27]), .B2(n1398), .ZN(n187) );
  AOI22_X1 U142 ( .A1(D[27]), .A2(n1416), .B1(C[27]), .B2(n1410), .ZN(n188) );
  NAND4_X1 U143 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U144 ( .A1(B[38]), .A2(n1405), .B1(A[38]), .B2(n1399), .ZN(n139) );
  AOI22_X1 U145 ( .A1(D[38]), .A2(n1417), .B1(C[38]), .B2(n1411), .ZN(n140) );
  AOI22_X1 U146 ( .A1(H[38]), .A2(n1441), .B1(G[38]), .B2(n1435), .ZN(n142) );
  NAND4_X1 U147 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U148 ( .A1(B[40]), .A2(n1405), .B1(A[40]), .B2(n1399), .ZN(n127) );
  AOI22_X1 U149 ( .A1(D[40]), .A2(n1417), .B1(C[40]), .B2(n1411), .ZN(n128) );
  AOI22_X1 U150 ( .A1(H[40]), .A2(n1441), .B1(G[40]), .B2(n1435), .ZN(n130) );
  NAND4_X1 U151 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U152 ( .A1(B[43]), .A2(n1406), .B1(A[43]), .B2(n1400), .ZN(n115) );
  AOI22_X1 U153 ( .A1(D[43]), .A2(n1418), .B1(C[43]), .B2(n1412), .ZN(n116) );
  AOI22_X1 U154 ( .A1(H[43]), .A2(n1442), .B1(G[43]), .B2(n1436), .ZN(n118) );
  NAND4_X1 U155 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U156 ( .A1(B[52]), .A2(n1406), .B1(A[52]), .B2(n1400), .ZN(n75) );
  AOI22_X1 U157 ( .A1(D[52]), .A2(n1418), .B1(C[52]), .B2(n1412), .ZN(n76) );
  AOI22_X1 U158 ( .A1(H[52]), .A2(n1442), .B1(G[52]), .B2(n1436), .ZN(n78) );
  NAND4_X1 U159 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U160 ( .A1(H[28]), .A2(n1440), .B1(G[28]), .B2(n1434), .ZN(n186) );
  AOI22_X1 U161 ( .A1(B[28]), .A2(n1404), .B1(A[28]), .B2(n1398), .ZN(n183) );
  AOI22_X1 U162 ( .A1(D[28]), .A2(n1416), .B1(C[28]), .B2(n1410), .ZN(n184) );
  NAND4_X1 U163 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U164 ( .A1(B[32]), .A2(n1405), .B1(A[32]), .B2(n1399), .ZN(n163) );
  AOI22_X1 U165 ( .A1(D[32]), .A2(n1417), .B1(C[32]), .B2(n1411), .ZN(n164) );
  AOI22_X1 U166 ( .A1(H[32]), .A2(n1441), .B1(G[32]), .B2(n1435), .ZN(n166) );
  NAND4_X1 U167 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U168 ( .A1(B[33]), .A2(n1405), .B1(A[33]), .B2(n1399), .ZN(n159) );
  AOI22_X1 U169 ( .A1(D[33]), .A2(n1417), .B1(C[33]), .B2(n1411), .ZN(n160) );
  AOI22_X1 U170 ( .A1(H[33]), .A2(n1441), .B1(G[33]), .B2(n1435), .ZN(n162) );
  NAND4_X1 U171 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U172 ( .A1(B[36]), .A2(n1405), .B1(A[36]), .B2(n1399), .ZN(n147) );
  AOI22_X1 U173 ( .A1(D[36]), .A2(n1417), .B1(C[36]), .B2(n1411), .ZN(n148) );
  AOI22_X1 U174 ( .A1(H[36]), .A2(n1441), .B1(G[36]), .B2(n1435), .ZN(n150) );
  NAND4_X1 U175 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U176 ( .A1(B[30]), .A2(n1404), .B1(A[30]), .B2(n1398), .ZN(n171) );
  AOI22_X1 U177 ( .A1(H[30]), .A2(n1440), .B1(G[30]), .B2(n1434), .ZN(n174) );
  AOI22_X1 U178 ( .A1(D[30]), .A2(n1416), .B1(C[30]), .B2(n1410), .ZN(n172) );
  NAND4_X1 U179 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U180 ( .A1(D[24]), .A2(n1416), .B1(C[24]), .B2(n1410), .ZN(n200) );
  AOI22_X1 U181 ( .A1(H[24]), .A2(n1440), .B1(G[24]), .B2(n1434), .ZN(n202) );
  AOI22_X1 U182 ( .A1(B[24]), .A2(n1404), .B1(A[24]), .B2(n1398), .ZN(n199) );
  NAND4_X1 U183 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U184 ( .A1(B[34]), .A2(n1405), .B1(A[34]), .B2(n1399), .ZN(n155) );
  AOI22_X1 U185 ( .A1(D[34]), .A2(n1417), .B1(C[34]), .B2(n1411), .ZN(n156) );
  AOI22_X1 U186 ( .A1(H[34]), .A2(n1441), .B1(G[34]), .B2(n1435), .ZN(n158) );
  NAND4_X1 U187 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U188 ( .A1(B[48]), .A2(n1406), .B1(A[48]), .B2(n1400), .ZN(n95) );
  AOI22_X1 U189 ( .A1(D[48]), .A2(n1418), .B1(C[48]), .B2(n1412), .ZN(n96) );
  AOI22_X1 U190 ( .A1(H[48]), .A2(n1442), .B1(G[48]), .B2(n1436), .ZN(n98) );
  NAND4_X1 U191 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U192 ( .A1(H[26]), .A2(n1440), .B1(G[26]), .B2(n1434), .ZN(n194) );
  AOI22_X1 U193 ( .A1(B[26]), .A2(n1404), .B1(A[26]), .B2(n1398), .ZN(n191) );
  AOI22_X1 U194 ( .A1(D[26]), .A2(n1416), .B1(C[26]), .B2(n1410), .ZN(n192) );
  NAND4_X1 U195 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U196 ( .A1(B[62]), .A2(n1407), .B1(A[62]), .B2(n1401), .ZN(n31) );
  AOI22_X1 U197 ( .A1(D[62]), .A2(n1419), .B1(C[62]), .B2(n1413), .ZN(n32) );
  AOI22_X1 U198 ( .A1(H[62]), .A2(n1443), .B1(G[62]), .B2(n1437), .ZN(n34) );
  NAND4_X1 U199 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U200 ( .A1(B[31]), .A2(n1405), .B1(A[31]), .B2(n1399), .ZN(n167) );
  AOI22_X1 U201 ( .A1(D[31]), .A2(n1417), .B1(C[31]), .B2(n1411), .ZN(n168) );
  AOI22_X1 U202 ( .A1(H[31]), .A2(n1441), .B1(G[31]), .B2(n1435), .ZN(n170) );
  NAND4_X1 U203 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U204 ( .A1(B[29]), .A2(n1404), .B1(A[29]), .B2(n1398), .ZN(n179) );
  AOI22_X1 U205 ( .A1(H[29]), .A2(n1440), .B1(G[29]), .B2(n1434), .ZN(n182) );
  AOI22_X1 U206 ( .A1(D[29]), .A2(n1416), .B1(C[29]), .B2(n1410), .ZN(n180) );
  NAND4_X1 U207 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U208 ( .A1(B[51]), .A2(n1406), .B1(A[51]), .B2(n1400), .ZN(n79) );
  AOI22_X1 U209 ( .A1(D[51]), .A2(n1418), .B1(C[51]), .B2(n1412), .ZN(n80) );
  AOI22_X1 U210 ( .A1(H[51]), .A2(n1442), .B1(G[51]), .B2(n1436), .ZN(n82) );
  NAND4_X1 U211 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U212 ( .A1(B[55]), .A2(n1407), .B1(A[55]), .B2(n1401), .ZN(n63) );
  AOI22_X1 U213 ( .A1(D[55]), .A2(n1419), .B1(C[55]), .B2(n1413), .ZN(n64) );
  AOI22_X1 U214 ( .A1(H[55]), .A2(n1443), .B1(G[55]), .B2(n1437), .ZN(n66) );
  NAND4_X1 U215 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U216 ( .A1(B[59]), .A2(n1407), .B1(A[59]), .B2(n1401), .ZN(n47) );
  AOI22_X1 U217 ( .A1(D[59]), .A2(n1419), .B1(C[59]), .B2(n1413), .ZN(n48) );
  AOI22_X1 U218 ( .A1(H[59]), .A2(n1443), .B1(G[59]), .B2(n1437), .ZN(n50) );
  AOI22_X1 U219 ( .A1(F[56]), .A2(n1431), .B1(E[56]), .B2(n1425), .ZN(n61) );
  AOI22_X1 U220 ( .A1(F[36]), .A2(n1429), .B1(E[36]), .B2(n1423), .ZN(n149) );
  AOI22_X1 U221 ( .A1(F[54]), .A2(n1431), .B1(E[54]), .B2(n1425), .ZN(n69) );
  AOI22_X1 U222 ( .A1(F[50]), .A2(n1430), .B1(E[50]), .B2(n1424), .ZN(n85) );
  AOI22_X1 U223 ( .A1(F[48]), .A2(n1430), .B1(E[48]), .B2(n1424), .ZN(n97) );
  AOI22_X1 U224 ( .A1(F[38]), .A2(n1429), .B1(E[38]), .B2(n1423), .ZN(n141) );
  NAND4_X1 U225 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U226 ( .A1(B[37]), .A2(n1405), .B1(A[37]), .B2(n1399), .ZN(n143) );
  AOI22_X1 U227 ( .A1(D[37]), .A2(n1417), .B1(C[37]), .B2(n1411), .ZN(n144) );
  AOI22_X1 U228 ( .A1(H[37]), .A2(n1441), .B1(G[37]), .B2(n1435), .ZN(n146) );
  NAND4_X1 U229 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U230 ( .A1(B[50]), .A2(n1406), .B1(A[50]), .B2(n1400), .ZN(n83) );
  AOI22_X1 U231 ( .A1(D[50]), .A2(n1418), .B1(C[50]), .B2(n1412), .ZN(n84) );
  AOI22_X1 U232 ( .A1(H[50]), .A2(n1442), .B1(G[50]), .B2(n1436), .ZN(n86) );
  NAND4_X1 U233 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U234 ( .A1(B[56]), .A2(n1407), .B1(A[56]), .B2(n1401), .ZN(n59) );
  AOI22_X1 U235 ( .A1(D[56]), .A2(n1419), .B1(C[56]), .B2(n1413), .ZN(n60) );
  AOI22_X1 U236 ( .A1(H[56]), .A2(n1443), .B1(G[56]), .B2(n1437), .ZN(n62) );
  NAND4_X1 U237 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U238 ( .A1(B[63]), .A2(n1407), .B1(A[63]), .B2(n1401), .ZN(n27) );
  AOI22_X1 U239 ( .A1(D[63]), .A2(n1419), .B1(C[63]), .B2(n1413), .ZN(n28) );
  AOI22_X1 U240 ( .A1(H[63]), .A2(n1443), .B1(G[63]), .B2(n1437), .ZN(n30) );
  AOI22_X1 U241 ( .A1(F[42]), .A2(n1430), .B1(E[42]), .B2(n1424), .ZN(n121) );
  AOI22_X1 U242 ( .A1(F[46]), .A2(n1430), .B1(E[46]), .B2(n1424), .ZN(n105) );
  NAND4_X1 U243 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U244 ( .A1(B[60]), .A2(n1407), .B1(A[60]), .B2(n1401), .ZN(n39) );
  AOI22_X1 U245 ( .A1(D[60]), .A2(n1419), .B1(C[60]), .B2(n1413), .ZN(n40) );
  AOI22_X1 U246 ( .A1(H[60]), .A2(n1443), .B1(G[60]), .B2(n1437), .ZN(n42) );
  NAND4_X1 U247 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U248 ( .A1(B[61]), .A2(n1407), .B1(A[61]), .B2(n1401), .ZN(n35) );
  AOI22_X1 U249 ( .A1(D[61]), .A2(n1419), .B1(C[61]), .B2(n1413), .ZN(n36) );
  AOI22_X1 U250 ( .A1(H[61]), .A2(n1443), .B1(G[61]), .B2(n1437), .ZN(n38) );
  NAND4_X1 U251 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U252 ( .A1(B[0]), .A2(n1403), .B1(A[0]), .B2(n1397), .ZN(n263) );
  AOI22_X1 U253 ( .A1(D[0]), .A2(n1415), .B1(C[0]), .B2(n1409), .ZN(n264) );
  AOI22_X1 U254 ( .A1(F[0]), .A2(n1427), .B1(E[0]), .B2(n1421), .ZN(n265) );
  AOI22_X1 U255 ( .A1(H[17]), .A2(n1439), .B1(G[17]), .B2(n1433), .ZN(n234) );
  AOI22_X1 U256 ( .A1(H[21]), .A2(n1440), .B1(G[21]), .B2(n1434), .ZN(n214) );
  AOI22_X1 U257 ( .A1(H[13]), .A2(n1439), .B1(G[13]), .B2(n1433), .ZN(n250) );
  AOI22_X1 U258 ( .A1(H[5]), .A2(n1443), .B1(G[5]), .B2(n1437), .ZN(n46) );
  AOI22_X1 U259 ( .A1(H[9]), .A2(n1444), .B1(G[9]), .B2(n1438), .ZN(n6) );
  AOI22_X1 U260 ( .A1(H[7]), .A2(n1444), .B1(G[7]), .B2(n1438), .ZN(n22) );
  AOI22_X1 U261 ( .A1(H[11]), .A2(n1439), .B1(G[11]), .B2(n1433), .ZN(n258) );
  AOI22_X1 U262 ( .A1(H[15]), .A2(n1439), .B1(G[15]), .B2(n1433), .ZN(n242) );
  AOI22_X1 U263 ( .A1(H[23]), .A2(n1440), .B1(G[23]), .B2(n1434), .ZN(n206) );
  AOI22_X1 U264 ( .A1(H[19]), .A2(n1439), .B1(G[19]), .B2(n1433), .ZN(n226) );
  AOI22_X1 U265 ( .A1(H[3]), .A2(n1441), .B1(G[3]), .B2(n1435), .ZN(n134) );
  AOI22_X1 U266 ( .A1(H[20]), .A2(n1440), .B1(G[20]), .B2(n1434), .ZN(n218) );
  AOI22_X1 U267 ( .A1(H[12]), .A2(n1439), .B1(G[12]), .B2(n1433), .ZN(n254) );
  AOI22_X1 U268 ( .A1(H[16]), .A2(n1439), .B1(G[16]), .B2(n1433), .ZN(n238) );
  AOI22_X1 U269 ( .A1(H[4]), .A2(n1442), .B1(G[4]), .B2(n1436), .ZN(n90) );
  AOI22_X1 U270 ( .A1(H[8]), .A2(n1444), .B1(G[8]), .B2(n1438), .ZN(n18) );
  AOI22_X1 U271 ( .A1(H[6]), .A2(n1444), .B1(G[6]), .B2(n1438), .ZN(n26) );
  AOI22_X1 U272 ( .A1(H[10]), .A2(n1439), .B1(G[10]), .B2(n1433), .ZN(n262) );
  AOI22_X1 U273 ( .A1(H[14]), .A2(n1439), .B1(G[14]), .B2(n1433), .ZN(n246) );
  AOI22_X1 U274 ( .A1(H[22]), .A2(n1440), .B1(G[22]), .B2(n1434), .ZN(n210) );
  AOI22_X1 U275 ( .A1(H[18]), .A2(n1439), .B1(G[18]), .B2(n1433), .ZN(n230) );
  AOI22_X1 U276 ( .A1(H[2]), .A2(n1440), .B1(G[2]), .B2(n1434), .ZN(n178) );
  AOI22_X1 U277 ( .A1(H[1]), .A2(n1439), .B1(G[1]), .B2(n1433), .ZN(n222) );
  NAND4_X1 U278 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U279 ( .A1(B[17]), .A2(n1403), .B1(A[17]), .B2(n1397), .ZN(n231) );
  AOI22_X1 U280 ( .A1(D[17]), .A2(n1415), .B1(C[17]), .B2(n1409), .ZN(n232) );
  AOI22_X1 U281 ( .A1(F[17]), .A2(n1427), .B1(E[17]), .B2(n1421), .ZN(n233) );
  NAND4_X1 U282 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U283 ( .A1(B[21]), .A2(n1404), .B1(A[21]), .B2(n1398), .ZN(n211) );
  AOI22_X1 U284 ( .A1(D[21]), .A2(n1416), .B1(C[21]), .B2(n1410), .ZN(n212) );
  AOI22_X1 U285 ( .A1(F[21]), .A2(n1428), .B1(E[21]), .B2(n1422), .ZN(n213) );
  NAND4_X1 U286 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U287 ( .A1(B[20]), .A2(n1404), .B1(A[20]), .B2(n1398), .ZN(n215) );
  AOI22_X1 U288 ( .A1(D[20]), .A2(n1416), .B1(C[20]), .B2(n1410), .ZN(n216) );
  AOI22_X1 U289 ( .A1(F[20]), .A2(n1428), .B1(E[20]), .B2(n1422), .ZN(n217) );
  NAND4_X1 U290 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U291 ( .A1(B[13]), .A2(n1403), .B1(A[13]), .B2(n1397), .ZN(n247) );
  AOI22_X1 U292 ( .A1(D[13]), .A2(n1415), .B1(C[13]), .B2(n1409), .ZN(n248) );
  AOI22_X1 U293 ( .A1(F[13]), .A2(n1427), .B1(E[13]), .B2(n1421), .ZN(n249) );
  NAND4_X1 U294 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U295 ( .A1(B[5]), .A2(n1407), .B1(A[5]), .B2(n1401), .ZN(n43) );
  AOI22_X1 U296 ( .A1(D[5]), .A2(n1419), .B1(C[5]), .B2(n1413), .ZN(n44) );
  AOI22_X1 U297 ( .A1(F[5]), .A2(n1431), .B1(E[5]), .B2(n1425), .ZN(n45) );
  NAND4_X1 U298 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U299 ( .A1(B[9]), .A2(n1408), .B1(A[9]), .B2(n1402), .ZN(n3) );
  AOI22_X1 U300 ( .A1(D[9]), .A2(n1420), .B1(C[9]), .B2(n1414), .ZN(n4) );
  AOI22_X1 U301 ( .A1(F[9]), .A2(n1432), .B1(E[9]), .B2(n1426), .ZN(n5) );
  NAND4_X1 U302 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U303 ( .A1(B[7]), .A2(n1408), .B1(A[7]), .B2(n1402), .ZN(n19) );
  AOI22_X1 U304 ( .A1(D[7]), .A2(n1420), .B1(C[7]), .B2(n1414), .ZN(n20) );
  AOI22_X1 U305 ( .A1(F[7]), .A2(n1432), .B1(E[7]), .B2(n1426), .ZN(n21) );
  NAND4_X1 U306 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U307 ( .A1(B[15]), .A2(n1403), .B1(A[15]), .B2(n1397), .ZN(n239) );
  AOI22_X1 U308 ( .A1(D[15]), .A2(n1415), .B1(C[15]), .B2(n1409), .ZN(n240) );
  AOI22_X1 U309 ( .A1(F[15]), .A2(n1427), .B1(E[15]), .B2(n1421), .ZN(n241) );
  NAND4_X1 U310 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U311 ( .A1(B[23]), .A2(n1404), .B1(A[23]), .B2(n1398), .ZN(n203) );
  AOI22_X1 U312 ( .A1(D[23]), .A2(n1416), .B1(C[23]), .B2(n1410), .ZN(n204) );
  AOI22_X1 U313 ( .A1(F[23]), .A2(n1428), .B1(E[23]), .B2(n1422), .ZN(n205) );
  NAND4_X1 U314 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U315 ( .A1(B[19]), .A2(n1403), .B1(A[19]), .B2(n1397), .ZN(n223) );
  AOI22_X1 U316 ( .A1(D[19]), .A2(n1415), .B1(C[19]), .B2(n1409), .ZN(n224) );
  AOI22_X1 U317 ( .A1(F[19]), .A2(n1427), .B1(E[19]), .B2(n1421), .ZN(n225) );
  NAND4_X1 U318 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U319 ( .A1(B[3]), .A2(n1405), .B1(A[3]), .B2(n1399), .ZN(n131) );
  AOI22_X1 U320 ( .A1(D[3]), .A2(n1417), .B1(C[3]), .B2(n1411), .ZN(n132) );
  AOI22_X1 U321 ( .A1(F[3]), .A2(n1429), .B1(E[3]), .B2(n1423), .ZN(n133) );
  NAND4_X1 U322 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U323 ( .A1(B[12]), .A2(n1403), .B1(A[12]), .B2(n1397), .ZN(n251) );
  AOI22_X1 U324 ( .A1(D[12]), .A2(n1415), .B1(C[12]), .B2(n1409), .ZN(n252) );
  AOI22_X1 U325 ( .A1(F[12]), .A2(n1427), .B1(E[12]), .B2(n1421), .ZN(n253) );
  NAND4_X1 U326 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U327 ( .A1(B[16]), .A2(n1403), .B1(A[16]), .B2(n1397), .ZN(n235) );
  AOI22_X1 U328 ( .A1(D[16]), .A2(n1415), .B1(C[16]), .B2(n1409), .ZN(n236) );
  AOI22_X1 U329 ( .A1(F[16]), .A2(n1427), .B1(E[16]), .B2(n1421), .ZN(n237) );
  NAND4_X1 U330 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U331 ( .A1(B[4]), .A2(n1406), .B1(A[4]), .B2(n1400), .ZN(n87) );
  AOI22_X1 U332 ( .A1(D[4]), .A2(n1418), .B1(C[4]), .B2(n1412), .ZN(n88) );
  AOI22_X1 U333 ( .A1(F[4]), .A2(n1430), .B1(E[4]), .B2(n1424), .ZN(n89) );
  NAND4_X1 U334 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U335 ( .A1(B[8]), .A2(n1408), .B1(A[8]), .B2(n1402), .ZN(n15) );
  AOI22_X1 U336 ( .A1(D[8]), .A2(n1420), .B1(C[8]), .B2(n1414), .ZN(n16) );
  AOI22_X1 U337 ( .A1(F[8]), .A2(n1432), .B1(E[8]), .B2(n1426), .ZN(n17) );
  NAND4_X1 U338 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U339 ( .A1(B[11]), .A2(n1403), .B1(A[11]), .B2(n1397), .ZN(n255) );
  AOI22_X1 U340 ( .A1(D[11]), .A2(n1415), .B1(C[11]), .B2(n1409), .ZN(n256) );
  AOI22_X1 U341 ( .A1(F[11]), .A2(n1427), .B1(E[11]), .B2(n1421), .ZN(n257) );
  NAND4_X1 U342 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U343 ( .A1(B[6]), .A2(n1408), .B1(A[6]), .B2(n1402), .ZN(n23) );
  AOI22_X1 U344 ( .A1(D[6]), .A2(n1420), .B1(C[6]), .B2(n1414), .ZN(n24) );
  AOI22_X1 U345 ( .A1(F[6]), .A2(n1432), .B1(E[6]), .B2(n1426), .ZN(n25) );
  NAND4_X1 U346 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U347 ( .A1(B[10]), .A2(n1403), .B1(A[10]), .B2(n1397), .ZN(n259) );
  AOI22_X1 U348 ( .A1(D[10]), .A2(n1415), .B1(C[10]), .B2(n1409), .ZN(n260) );
  AOI22_X1 U349 ( .A1(F[10]), .A2(n1427), .B1(E[10]), .B2(n1421), .ZN(n261) );
  NAND4_X1 U350 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U351 ( .A1(B[14]), .A2(n1403), .B1(A[14]), .B2(n1397), .ZN(n243) );
  AOI22_X1 U352 ( .A1(D[14]), .A2(n1415), .B1(C[14]), .B2(n1409), .ZN(n244) );
  AOI22_X1 U353 ( .A1(F[14]), .A2(n1427), .B1(E[14]), .B2(n1421), .ZN(n245) );
  NAND4_X1 U354 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U355 ( .A1(B[22]), .A2(n1404), .B1(A[22]), .B2(n1398), .ZN(n207) );
  AOI22_X1 U356 ( .A1(D[22]), .A2(n1416), .B1(C[22]), .B2(n1410), .ZN(n208) );
  AOI22_X1 U357 ( .A1(F[22]), .A2(n1428), .B1(E[22]), .B2(n1422), .ZN(n209) );
  NAND4_X1 U358 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U359 ( .A1(B[18]), .A2(n1403), .B1(A[18]), .B2(n1397), .ZN(n227) );
  AOI22_X1 U360 ( .A1(D[18]), .A2(n1415), .B1(C[18]), .B2(n1409), .ZN(n228) );
  AOI22_X1 U361 ( .A1(F[18]), .A2(n1427), .B1(E[18]), .B2(n1421), .ZN(n229) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1404), .B1(A[2]), .B2(n1398), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1416), .B1(C[2]), .B2(n1410), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1428), .B1(E[2]), .B2(n1422), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1403), .B1(A[1]), .B2(n1397), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1415), .B1(C[1]), .B2(n1409), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1427), .B1(E[1]), .B2(n1421), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1439), .B1(G[0]), .B2(n1433), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1402) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1408) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1414) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1420) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1426) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1432) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1438) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1444) );
endmodule


module MUX81_GENERIC_NBIT64_3 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442;

  BUF_X1 U1 ( .A(n13), .Z(n1402) );
  BUF_X1 U2 ( .A(n13), .Z(n1400) );
  BUF_X1 U3 ( .A(n13), .Z(n1401) );
  BUF_X1 U4 ( .A(n12), .Z(n1408) );
  BUF_X1 U5 ( .A(n12), .Z(n1406) );
  BUF_X1 U6 ( .A(n12), .Z(n1407) );
  BUF_X1 U7 ( .A(n8), .Z(n1431) );
  BUF_X1 U8 ( .A(n8), .Z(n1430) );
  BUF_X1 U9 ( .A(n10), .Z(n1420) );
  BUF_X1 U10 ( .A(n8), .Z(n1432) );
  BUF_X1 U11 ( .A(n10), .Z(n1418) );
  BUF_X1 U12 ( .A(n10), .Z(n1419) );
  BUF_X1 U13 ( .A(n13), .Z(n1403) );
  BUF_X1 U14 ( .A(n12), .Z(n1409) );
  BUF_X1 U15 ( .A(n10), .Z(n1421) );
  BUF_X1 U16 ( .A(n8), .Z(n1433) );
  BUF_X1 U17 ( .A(n11), .Z(n1414) );
  BUF_X1 U18 ( .A(n11), .Z(n1412) );
  BUF_X1 U19 ( .A(n11), .Z(n1413) );
  BUF_X1 U20 ( .A(n11), .Z(n1411) );
  BUF_X1 U21 ( .A(n13), .Z(n1399) );
  BUF_X1 U22 ( .A(n11), .Z(n1415) );
  BUF_X1 U23 ( .A(n7), .Z(n1435) );
  BUF_X1 U24 ( .A(n7), .Z(n1437) );
  BUF_X1 U25 ( .A(n7), .Z(n1436) );
  BUF_X1 U26 ( .A(n9), .Z(n1426) );
  BUF_X1 U27 ( .A(n7), .Z(n1438) );
  BUF_X1 U28 ( .A(n9), .Z(n1427) );
  BUF_X1 U29 ( .A(n9), .Z(n1424) );
  BUF_X1 U30 ( .A(n9), .Z(n1425) );
  BUF_X1 U31 ( .A(n9), .Z(n1423) );
  BUF_X1 U32 ( .A(n7), .Z(n1439) );
  BUF_X1 U33 ( .A(n14), .Z(n1396) );
  BUF_X1 U34 ( .A(n14), .Z(n1394) );
  BUF_X1 U35 ( .A(n14), .Z(n1395) );
  BUF_X1 U36 ( .A(n12), .Z(n1405) );
  BUF_X1 U37 ( .A(n14), .Z(n1393) );
  BUF_X1 U38 ( .A(n14), .Z(n1397) );
  BUF_X1 U39 ( .A(n8), .Z(n1429) );
  BUF_X1 U40 ( .A(n10), .Z(n1417) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1441), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1442), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1442), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1442), .A2(n1441), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1441) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1442) );
  NOR3_X1 U47 ( .A1(n1442), .A2(SEL[2]), .A3(n1441), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1441), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U52 ( .A1(B[52]), .A2(n1402), .B1(A[52]), .B2(n1396), .ZN(n75) );
  AOI22_X1 U53 ( .A1(D[52]), .A2(n1414), .B1(C[52]), .B2(n1408), .ZN(n76) );
  AOI22_X1 U54 ( .A1(H[52]), .A2(n1438), .B1(G[52]), .B2(n1432), .ZN(n78) );
  AOI22_X1 U55 ( .A1(F[62]), .A2(n1427), .B1(E[62]), .B2(n1421), .ZN(n33) );
  AOI22_X1 U56 ( .A1(F[55]), .A2(n1427), .B1(E[55]), .B2(n1421), .ZN(n65) );
  AOI22_X1 U57 ( .A1(F[61]), .A2(n1427), .B1(E[61]), .B2(n1421), .ZN(n37) );
  NAND4_X1 U58 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U59 ( .A1(B[48]), .A2(n1402), .B1(A[48]), .B2(n1396), .ZN(n95) );
  AOI22_X1 U60 ( .A1(D[48]), .A2(n1414), .B1(C[48]), .B2(n1408), .ZN(n96) );
  AOI22_X1 U61 ( .A1(H[48]), .A2(n1438), .B1(G[48]), .B2(n1432), .ZN(n98) );
  NAND4_X1 U62 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U63 ( .A1(B[45]), .A2(n1402), .B1(A[45]), .B2(n1396), .ZN(n107) );
  AOI22_X1 U64 ( .A1(D[45]), .A2(n1414), .B1(C[45]), .B2(n1408), .ZN(n108) );
  AOI22_X1 U65 ( .A1(H[45]), .A2(n1438), .B1(G[45]), .B2(n1432), .ZN(n110) );
  NAND4_X1 U66 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U67 ( .A1(B[54]), .A2(n1403), .B1(A[54]), .B2(n1397), .ZN(n67) );
  AOI22_X1 U68 ( .A1(D[54]), .A2(n1415), .B1(C[54]), .B2(n1409), .ZN(n68) );
  AOI22_X1 U69 ( .A1(H[54]), .A2(n1439), .B1(G[54]), .B2(n1433), .ZN(n70) );
  NAND4_X1 U70 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U71 ( .A1(B[56]), .A2(n1403), .B1(A[56]), .B2(n1397), .ZN(n59) );
  AOI22_X1 U72 ( .A1(D[56]), .A2(n1415), .B1(C[56]), .B2(n1409), .ZN(n60) );
  AOI22_X1 U73 ( .A1(H[56]), .A2(n1439), .B1(G[56]), .B2(n1433), .ZN(n62) );
  NAND4_X1 U74 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U75 ( .A1(B[46]), .A2(n1402), .B1(A[46]), .B2(n1396), .ZN(n103) );
  AOI22_X1 U76 ( .A1(D[46]), .A2(n1414), .B1(C[46]), .B2(n1408), .ZN(n104) );
  AOI22_X1 U77 ( .A1(H[46]), .A2(n1438), .B1(G[46]), .B2(n1432), .ZN(n106) );
  NAND4_X1 U78 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U79 ( .A1(B[55]), .A2(n1403), .B1(A[55]), .B2(n1397), .ZN(n63) );
  AOI22_X1 U80 ( .A1(D[55]), .A2(n1415), .B1(C[55]), .B2(n1409), .ZN(n64) );
  AOI22_X1 U81 ( .A1(H[55]), .A2(n1439), .B1(G[55]), .B2(n1433), .ZN(n66) );
  AOI22_X1 U82 ( .A1(F[45]), .A2(n1426), .B1(E[45]), .B2(n1420), .ZN(n109) );
  AOI22_X1 U83 ( .A1(F[47]), .A2(n1426), .B1(E[47]), .B2(n1420), .ZN(n101) );
  AOI22_X1 U84 ( .A1(F[49]), .A2(n1426), .B1(E[49]), .B2(n1420), .ZN(n93) );
  AOI22_X1 U85 ( .A1(F[48]), .A2(n1426), .B1(E[48]), .B2(n1420), .ZN(n97) );
  AOI22_X1 U86 ( .A1(F[53]), .A2(n1427), .B1(E[53]), .B2(n1421), .ZN(n73) );
  AOI22_X1 U87 ( .A1(F[51]), .A2(n1426), .B1(E[51]), .B2(n1420), .ZN(n81) );
  AOI22_X1 U88 ( .A1(F[57]), .A2(n1427), .B1(E[57]), .B2(n1421), .ZN(n57) );
  AOI22_X1 U89 ( .A1(F[59]), .A2(n1427), .B1(E[59]), .B2(n1421), .ZN(n49) );
  AOI22_X1 U90 ( .A1(F[58]), .A2(n1427), .B1(E[58]), .B2(n1421), .ZN(n53) );
  AOI22_X1 U91 ( .A1(F[63]), .A2(n1427), .B1(E[63]), .B2(n1421), .ZN(n29) );
  NAND4_X1 U92 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U93 ( .A1(B[50]), .A2(n1402), .B1(A[50]), .B2(n1396), .ZN(n83) );
  AOI22_X1 U94 ( .A1(D[50]), .A2(n1414), .B1(C[50]), .B2(n1408), .ZN(n84) );
  AOI22_X1 U95 ( .A1(H[50]), .A2(n1438), .B1(G[50]), .B2(n1432), .ZN(n86) );
  NAND4_X1 U96 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U97 ( .A1(B[53]), .A2(n1403), .B1(A[53]), .B2(n1397), .ZN(n71) );
  AOI22_X1 U98 ( .A1(D[53]), .A2(n1415), .B1(C[53]), .B2(n1409), .ZN(n72) );
  AOI22_X1 U99 ( .A1(H[53]), .A2(n1439), .B1(G[53]), .B2(n1433), .ZN(n74) );
  NAND4_X1 U100 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U101 ( .A1(B[59]), .A2(n1403), .B1(A[59]), .B2(n1397), .ZN(n47) );
  AOI22_X1 U102 ( .A1(D[59]), .A2(n1415), .B1(C[59]), .B2(n1409), .ZN(n48) );
  AOI22_X1 U103 ( .A1(H[59]), .A2(n1439), .B1(G[59]), .B2(n1433), .ZN(n50) );
  NAND4_X1 U104 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U105 ( .A1(B[49]), .A2(n1402), .B1(A[49]), .B2(n1396), .ZN(n91) );
  AOI22_X1 U106 ( .A1(D[49]), .A2(n1414), .B1(C[49]), .B2(n1408), .ZN(n92) );
  AOI22_X1 U107 ( .A1(H[49]), .A2(n1438), .B1(G[49]), .B2(n1432), .ZN(n94) );
  NAND4_X1 U108 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U109 ( .A1(B[47]), .A2(n1402), .B1(A[47]), .B2(n1396), .ZN(n99) );
  AOI22_X1 U110 ( .A1(D[47]), .A2(n1414), .B1(C[47]), .B2(n1408), .ZN(n100) );
  AOI22_X1 U111 ( .A1(H[47]), .A2(n1438), .B1(G[47]), .B2(n1432), .ZN(n102) );
  AOI22_X1 U112 ( .A1(F[60]), .A2(n1427), .B1(E[60]), .B2(n1421), .ZN(n41) );
  AOI22_X1 U113 ( .A1(F[56]), .A2(n1427), .B1(E[56]), .B2(n1421), .ZN(n61) );
  AOI22_X1 U114 ( .A1(F[52]), .A2(n1426), .B1(E[52]), .B2(n1420), .ZN(n77) );
  AOI22_X1 U115 ( .A1(F[46]), .A2(n1426), .B1(E[46]), .B2(n1420), .ZN(n105) );
  NAND4_X1 U116 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U117 ( .A1(B[60]), .A2(n1403), .B1(A[60]), .B2(n1397), .ZN(n39) );
  AOI22_X1 U118 ( .A1(D[60]), .A2(n1415), .B1(C[60]), .B2(n1409), .ZN(n40) );
  AOI22_X1 U119 ( .A1(H[60]), .A2(n1439), .B1(G[60]), .B2(n1433), .ZN(n42) );
  NAND4_X1 U120 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U121 ( .A1(B[57]), .A2(n1403), .B1(A[57]), .B2(n1397), .ZN(n55) );
  AOI22_X1 U122 ( .A1(D[57]), .A2(n1415), .B1(C[57]), .B2(n1409), .ZN(n56) );
  AOI22_X1 U123 ( .A1(H[57]), .A2(n1439), .B1(G[57]), .B2(n1433), .ZN(n58) );
  NAND4_X1 U124 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U125 ( .A1(B[51]), .A2(n1402), .B1(A[51]), .B2(n1396), .ZN(n79) );
  AOI22_X1 U126 ( .A1(D[51]), .A2(n1414), .B1(C[51]), .B2(n1408), .ZN(n80) );
  AOI22_X1 U127 ( .A1(H[51]), .A2(n1438), .B1(G[51]), .B2(n1432), .ZN(n82) );
  NAND4_X1 U128 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U129 ( .A1(B[61]), .A2(n1403), .B1(A[61]), .B2(n1397), .ZN(n35) );
  AOI22_X1 U130 ( .A1(D[61]), .A2(n1415), .B1(C[61]), .B2(n1409), .ZN(n36) );
  AOI22_X1 U131 ( .A1(H[61]), .A2(n1439), .B1(G[61]), .B2(n1433), .ZN(n38) );
  NAND4_X1 U132 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U133 ( .A1(B[62]), .A2(n1403), .B1(A[62]), .B2(n1397), .ZN(n31) );
  AOI22_X1 U134 ( .A1(D[62]), .A2(n1415), .B1(C[62]), .B2(n1409), .ZN(n32) );
  AOI22_X1 U135 ( .A1(H[62]), .A2(n1439), .B1(G[62]), .B2(n1433), .ZN(n34) );
  AOI22_X1 U136 ( .A1(F[50]), .A2(n1426), .B1(E[50]), .B2(n1420), .ZN(n85) );
  NAND4_X1 U137 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U138 ( .A1(B[58]), .A2(n1403), .B1(A[58]), .B2(n1397), .ZN(n51) );
  AOI22_X1 U139 ( .A1(D[58]), .A2(n1415), .B1(C[58]), .B2(n1409), .ZN(n52) );
  AOI22_X1 U140 ( .A1(H[58]), .A2(n1439), .B1(G[58]), .B2(n1433), .ZN(n54) );
  NAND4_X1 U141 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U142 ( .A1(B[63]), .A2(n1403), .B1(A[63]), .B2(n1397), .ZN(n27) );
  AOI22_X1 U143 ( .A1(D[63]), .A2(n1415), .B1(C[63]), .B2(n1409), .ZN(n28) );
  AOI22_X1 U144 ( .A1(H[63]), .A2(n1439), .B1(G[63]), .B2(n1433), .ZN(n30) );
  AOI22_X1 U145 ( .A1(F[54]), .A2(n1427), .B1(E[54]), .B2(n1421), .ZN(n69) );
  AOI22_X1 U146 ( .A1(F[35]), .A2(n1425), .B1(E[35]), .B2(n1419), .ZN(n153) );
  AOI22_X1 U147 ( .A1(F[31]), .A2(n1425), .B1(E[31]), .B2(n1419), .ZN(n169) );
  AOI22_X1 U148 ( .A1(F[33]), .A2(n1425), .B1(E[33]), .B2(n1419), .ZN(n161) );
  AOI22_X1 U149 ( .A1(F[29]), .A2(n1424), .B1(E[29]), .B2(n1418), .ZN(n181) );
  AOI22_X1 U150 ( .A1(F[39]), .A2(n1425), .B1(E[39]), .B2(n1419), .ZN(n137) );
  AOI22_X1 U151 ( .A1(F[37]), .A2(n1425), .B1(E[37]), .B2(n1419), .ZN(n145) );
  AOI22_X1 U152 ( .A1(F[41]), .A2(n1425), .B1(E[41]), .B2(n1419), .ZN(n125) );
  AOI22_X1 U153 ( .A1(F[38]), .A2(n1425), .B1(E[38]), .B2(n1419), .ZN(n141) );
  AOI22_X1 U154 ( .A1(F[43]), .A2(n1426), .B1(E[43]), .B2(n1420), .ZN(n117) );
  AOI22_X1 U155 ( .A1(F[34]), .A2(n1425), .B1(E[34]), .B2(n1419), .ZN(n157) );
  AOI22_X1 U156 ( .A1(F[26]), .A2(n1424), .B1(E[26]), .B2(n1418), .ZN(n193) );
  AOI22_X1 U157 ( .A1(D[28]), .A2(n1412), .B1(C[28]), .B2(n1406), .ZN(n184) );
  AOI22_X1 U158 ( .A1(D[30]), .A2(n1412), .B1(C[30]), .B2(n1406), .ZN(n172) );
  AOI22_X1 U159 ( .A1(D[27]), .A2(n1412), .B1(C[27]), .B2(n1406), .ZN(n188) );
  NAND4_X1 U160 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U161 ( .A1(B[35]), .A2(n1401), .B1(A[35]), .B2(n1395), .ZN(n151) );
  AOI22_X1 U162 ( .A1(D[35]), .A2(n1413), .B1(C[35]), .B2(n1407), .ZN(n152) );
  AOI22_X1 U163 ( .A1(H[35]), .A2(n1437), .B1(G[35]), .B2(n1431), .ZN(n154) );
  NAND4_X1 U164 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U165 ( .A1(B[40]), .A2(n1401), .B1(A[40]), .B2(n1395), .ZN(n127) );
  AOI22_X1 U166 ( .A1(D[40]), .A2(n1413), .B1(C[40]), .B2(n1407), .ZN(n128) );
  AOI22_X1 U167 ( .A1(H[40]), .A2(n1437), .B1(G[40]), .B2(n1431), .ZN(n130) );
  NAND4_X1 U168 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U169 ( .A1(B[42]), .A2(n1402), .B1(A[42]), .B2(n1396), .ZN(n119) );
  AOI22_X1 U170 ( .A1(D[42]), .A2(n1414), .B1(C[42]), .B2(n1408), .ZN(n120) );
  AOI22_X1 U171 ( .A1(H[42]), .A2(n1438), .B1(G[42]), .B2(n1432), .ZN(n122) );
  NAND4_X1 U172 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U173 ( .A1(H[27]), .A2(n1436), .B1(G[27]), .B2(n1430), .ZN(n190) );
  AOI22_X1 U174 ( .A1(B[27]), .A2(n1400), .B1(A[27]), .B2(n1394), .ZN(n187) );
  AOI22_X1 U175 ( .A1(F[27]), .A2(n1424), .B1(E[27]), .B2(n1418), .ZN(n189) );
  NAND4_X1 U176 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U177 ( .A1(B[33]), .A2(n1401), .B1(A[33]), .B2(n1395), .ZN(n159) );
  AOI22_X1 U178 ( .A1(H[33]), .A2(n1437), .B1(G[33]), .B2(n1431), .ZN(n162) );
  AOI22_X1 U179 ( .A1(D[33]), .A2(n1413), .B1(C[33]), .B2(n1407), .ZN(n160) );
  NAND4_X1 U180 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U181 ( .A1(H[32]), .A2(n1437), .B1(G[32]), .B2(n1431), .ZN(n166) );
  AOI22_X1 U182 ( .A1(B[32]), .A2(n1401), .B1(A[32]), .B2(n1395), .ZN(n163) );
  AOI22_X1 U183 ( .A1(D[32]), .A2(n1413), .B1(C[32]), .B2(n1407), .ZN(n164) );
  NAND4_X1 U184 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U185 ( .A1(B[39]), .A2(n1401), .B1(A[39]), .B2(n1395), .ZN(n135) );
  AOI22_X1 U186 ( .A1(D[39]), .A2(n1413), .B1(C[39]), .B2(n1407), .ZN(n136) );
  AOI22_X1 U187 ( .A1(H[39]), .A2(n1437), .B1(G[39]), .B2(n1431), .ZN(n138) );
  NAND4_X1 U188 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U189 ( .A1(B[36]), .A2(n1401), .B1(A[36]), .B2(n1395), .ZN(n147) );
  AOI22_X1 U190 ( .A1(D[36]), .A2(n1413), .B1(C[36]), .B2(n1407), .ZN(n148) );
  AOI22_X1 U191 ( .A1(H[36]), .A2(n1437), .B1(G[36]), .B2(n1431), .ZN(n150) );
  NAND4_X1 U192 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U193 ( .A1(B[37]), .A2(n1401), .B1(A[37]), .B2(n1395), .ZN(n143) );
  AOI22_X1 U194 ( .A1(D[37]), .A2(n1413), .B1(C[37]), .B2(n1407), .ZN(n144) );
  AOI22_X1 U195 ( .A1(H[37]), .A2(n1437), .B1(G[37]), .B2(n1431), .ZN(n146) );
  NAND4_X1 U196 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U197 ( .A1(H[28]), .A2(n1436), .B1(G[28]), .B2(n1430), .ZN(n186) );
  AOI22_X1 U198 ( .A1(B[28]), .A2(n1400), .B1(A[28]), .B2(n1394), .ZN(n183) );
  AOI22_X1 U199 ( .A1(F[28]), .A2(n1424), .B1(E[28]), .B2(n1418), .ZN(n185) );
  NAND4_X1 U200 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U201 ( .A1(B[38]), .A2(n1401), .B1(A[38]), .B2(n1395), .ZN(n139) );
  AOI22_X1 U202 ( .A1(D[38]), .A2(n1413), .B1(C[38]), .B2(n1407), .ZN(n140) );
  AOI22_X1 U203 ( .A1(H[38]), .A2(n1437), .B1(G[38]), .B2(n1431), .ZN(n142) );
  NAND4_X1 U204 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U205 ( .A1(H[30]), .A2(n1436), .B1(G[30]), .B2(n1430), .ZN(n174) );
  AOI22_X1 U206 ( .A1(B[30]), .A2(n1400), .B1(A[30]), .B2(n1394), .ZN(n171) );
  AOI22_X1 U207 ( .A1(F[30]), .A2(n1424), .B1(E[30]), .B2(n1418), .ZN(n173) );
  NAND4_X1 U208 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U209 ( .A1(B[44]), .A2(n1402), .B1(A[44]), .B2(n1396), .ZN(n111) );
  AOI22_X1 U210 ( .A1(D[44]), .A2(n1414), .B1(C[44]), .B2(n1408), .ZN(n112) );
  AOI22_X1 U211 ( .A1(H[44]), .A2(n1438), .B1(G[44]), .B2(n1432), .ZN(n114) );
  NAND4_X1 U212 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U213 ( .A1(B[34]), .A2(n1401), .B1(A[34]), .B2(n1395), .ZN(n155) );
  AOI22_X1 U214 ( .A1(H[34]), .A2(n1437), .B1(G[34]), .B2(n1431), .ZN(n158) );
  AOI22_X1 U215 ( .A1(D[34]), .A2(n1413), .B1(C[34]), .B2(n1407), .ZN(n156) );
  NAND4_X1 U216 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U217 ( .A1(D[26]), .A2(n1412), .B1(C[26]), .B2(n1406), .ZN(n192) );
  AOI22_X1 U218 ( .A1(H[26]), .A2(n1436), .B1(G[26]), .B2(n1430), .ZN(n194) );
  AOI22_X1 U219 ( .A1(B[26]), .A2(n1400), .B1(A[26]), .B2(n1394), .ZN(n191) );
  NAND4_X1 U220 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U221 ( .A1(H[29]), .A2(n1436), .B1(G[29]), .B2(n1430), .ZN(n182) );
  AOI22_X1 U222 ( .A1(B[29]), .A2(n1400), .B1(A[29]), .B2(n1394), .ZN(n179) );
  AOI22_X1 U223 ( .A1(D[29]), .A2(n1412), .B1(C[29]), .B2(n1406), .ZN(n180) );
  NAND4_X1 U224 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U225 ( .A1(H[31]), .A2(n1437), .B1(G[31]), .B2(n1431), .ZN(n170) );
  AOI22_X1 U226 ( .A1(B[31]), .A2(n1401), .B1(A[31]), .B2(n1395), .ZN(n167) );
  AOI22_X1 U227 ( .A1(D[31]), .A2(n1413), .B1(C[31]), .B2(n1407), .ZN(n168) );
  NAND4_X1 U228 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U229 ( .A1(B[41]), .A2(n1401), .B1(A[41]), .B2(n1395), .ZN(n123) );
  AOI22_X1 U230 ( .A1(D[41]), .A2(n1413), .B1(C[41]), .B2(n1407), .ZN(n124) );
  AOI22_X1 U231 ( .A1(H[41]), .A2(n1437), .B1(G[41]), .B2(n1431), .ZN(n126) );
  AOI22_X1 U232 ( .A1(F[44]), .A2(n1426), .B1(E[44]), .B2(n1420), .ZN(n113) );
  AOI22_X1 U233 ( .A1(F[36]), .A2(n1425), .B1(E[36]), .B2(n1419), .ZN(n149) );
  AOI22_X1 U234 ( .A1(F[32]), .A2(n1425), .B1(E[32]), .B2(n1419), .ZN(n165) );
  AOI22_X1 U235 ( .A1(F[40]), .A2(n1425), .B1(E[40]), .B2(n1419), .ZN(n129) );
  AOI22_X1 U236 ( .A1(F[42]), .A2(n1426), .B1(E[42]), .B2(n1420), .ZN(n121) );
  NAND4_X1 U237 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U238 ( .A1(B[43]), .A2(n1402), .B1(A[43]), .B2(n1396), .ZN(n115) );
  AOI22_X1 U239 ( .A1(D[43]), .A2(n1414), .B1(C[43]), .B2(n1408), .ZN(n116) );
  AOI22_X1 U240 ( .A1(H[43]), .A2(n1438), .B1(G[43]), .B2(n1432), .ZN(n118) );
  NAND4_X1 U241 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U242 ( .A1(B[0]), .A2(n1399), .B1(A[0]), .B2(n1393), .ZN(n263) );
  AOI22_X1 U243 ( .A1(D[0]), .A2(n1411), .B1(C[0]), .B2(n1405), .ZN(n264) );
  AOI22_X1 U244 ( .A1(F[0]), .A2(n1423), .B1(E[0]), .B2(n1417), .ZN(n265) );
  AOI22_X1 U245 ( .A1(H[17]), .A2(n1435), .B1(G[17]), .B2(n1429), .ZN(n234) );
  AOI22_X1 U246 ( .A1(H[21]), .A2(n1436), .B1(G[21]), .B2(n1430), .ZN(n214) );
  AOI22_X1 U247 ( .A1(H[13]), .A2(n1435), .B1(G[13]), .B2(n1429), .ZN(n250) );
  AOI22_X1 U248 ( .A1(H[25]), .A2(n1436), .B1(G[25]), .B2(n1430), .ZN(n198) );
  AOI22_X1 U249 ( .A1(H[5]), .A2(n1439), .B1(G[5]), .B2(n1433), .ZN(n46) );
  AOI22_X1 U250 ( .A1(H[9]), .A2(n1440), .B1(G[9]), .B2(n1434), .ZN(n6) );
  AOI22_X1 U251 ( .A1(H[7]), .A2(n1440), .B1(G[7]), .B2(n1434), .ZN(n22) );
  AOI22_X1 U252 ( .A1(H[11]), .A2(n1435), .B1(G[11]), .B2(n1429), .ZN(n258) );
  AOI22_X1 U253 ( .A1(H[15]), .A2(n1435), .B1(G[15]), .B2(n1429), .ZN(n242) );
  AOI22_X1 U254 ( .A1(H[23]), .A2(n1436), .B1(G[23]), .B2(n1430), .ZN(n206) );
  AOI22_X1 U255 ( .A1(H[19]), .A2(n1435), .B1(G[19]), .B2(n1429), .ZN(n226) );
  AOI22_X1 U256 ( .A1(H[3]), .A2(n1437), .B1(G[3]), .B2(n1431), .ZN(n134) );
  AOI22_X1 U257 ( .A1(H[20]), .A2(n1436), .B1(G[20]), .B2(n1430), .ZN(n218) );
  AOI22_X1 U258 ( .A1(H[12]), .A2(n1435), .B1(G[12]), .B2(n1429), .ZN(n254) );
  AOI22_X1 U259 ( .A1(H[16]), .A2(n1435), .B1(G[16]), .B2(n1429), .ZN(n238) );
  AOI22_X1 U260 ( .A1(H[24]), .A2(n1436), .B1(G[24]), .B2(n1430), .ZN(n202) );
  AOI22_X1 U261 ( .A1(H[4]), .A2(n1438), .B1(G[4]), .B2(n1432), .ZN(n90) );
  AOI22_X1 U262 ( .A1(H[8]), .A2(n1440), .B1(G[8]), .B2(n1434), .ZN(n18) );
  AOI22_X1 U263 ( .A1(H[6]), .A2(n1440), .B1(G[6]), .B2(n1434), .ZN(n26) );
  AOI22_X1 U264 ( .A1(H[10]), .A2(n1435), .B1(G[10]), .B2(n1429), .ZN(n262) );
  AOI22_X1 U265 ( .A1(H[14]), .A2(n1435), .B1(G[14]), .B2(n1429), .ZN(n246) );
  AOI22_X1 U266 ( .A1(H[22]), .A2(n1436), .B1(G[22]), .B2(n1430), .ZN(n210) );
  AOI22_X1 U267 ( .A1(H[18]), .A2(n1435), .B1(G[18]), .B2(n1429), .ZN(n230) );
  AOI22_X1 U268 ( .A1(H[2]), .A2(n1436), .B1(G[2]), .B2(n1430), .ZN(n178) );
  AOI22_X1 U269 ( .A1(H[1]), .A2(n1435), .B1(G[1]), .B2(n1429), .ZN(n222) );
  NAND4_X1 U270 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U271 ( .A1(B[17]), .A2(n1399), .B1(A[17]), .B2(n1393), .ZN(n231) );
  AOI22_X1 U272 ( .A1(D[17]), .A2(n1411), .B1(C[17]), .B2(n1405), .ZN(n232) );
  AOI22_X1 U273 ( .A1(F[17]), .A2(n1423), .B1(E[17]), .B2(n1417), .ZN(n233) );
  NAND4_X1 U274 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U275 ( .A1(B[21]), .A2(n1400), .B1(A[21]), .B2(n1394), .ZN(n211) );
  AOI22_X1 U276 ( .A1(D[21]), .A2(n1412), .B1(C[21]), .B2(n1406), .ZN(n212) );
  AOI22_X1 U277 ( .A1(F[21]), .A2(n1424), .B1(E[21]), .B2(n1418), .ZN(n213) );
  NAND4_X1 U278 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U279 ( .A1(B[20]), .A2(n1400), .B1(A[20]), .B2(n1394), .ZN(n215) );
  AOI22_X1 U280 ( .A1(D[20]), .A2(n1412), .B1(C[20]), .B2(n1406), .ZN(n216) );
  AOI22_X1 U281 ( .A1(F[20]), .A2(n1424), .B1(E[20]), .B2(n1418), .ZN(n217) );
  NAND4_X1 U282 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U283 ( .A1(B[13]), .A2(n1399), .B1(A[13]), .B2(n1393), .ZN(n247) );
  AOI22_X1 U284 ( .A1(D[13]), .A2(n1411), .B1(C[13]), .B2(n1405), .ZN(n248) );
  AOI22_X1 U285 ( .A1(F[13]), .A2(n1423), .B1(E[13]), .B2(n1417), .ZN(n249) );
  NAND4_X1 U286 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U287 ( .A1(B[16]), .A2(n1399), .B1(A[16]), .B2(n1393), .ZN(n235) );
  AOI22_X1 U288 ( .A1(D[16]), .A2(n1411), .B1(C[16]), .B2(n1405), .ZN(n236) );
  AOI22_X1 U289 ( .A1(F[16]), .A2(n1423), .B1(E[16]), .B2(n1417), .ZN(n237) );
  NAND4_X1 U290 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U291 ( .A1(B[24]), .A2(n1400), .B1(A[24]), .B2(n1394), .ZN(n199) );
  AOI22_X1 U292 ( .A1(D[24]), .A2(n1412), .B1(C[24]), .B2(n1406), .ZN(n200) );
  AOI22_X1 U293 ( .A1(F[24]), .A2(n1424), .B1(E[24]), .B2(n1418), .ZN(n201) );
  NAND4_X1 U294 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U295 ( .A1(B[25]), .A2(n1400), .B1(A[25]), .B2(n1394), .ZN(n195) );
  AOI22_X1 U296 ( .A1(D[25]), .A2(n1412), .B1(C[25]), .B2(n1406), .ZN(n196) );
  AOI22_X1 U297 ( .A1(F[25]), .A2(n1424), .B1(E[25]), .B2(n1418), .ZN(n197) );
  NAND4_X1 U298 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U299 ( .A1(B[8]), .A2(n1404), .B1(A[8]), .B2(n1398), .ZN(n15) );
  AOI22_X1 U300 ( .A1(D[8]), .A2(n1416), .B1(C[8]), .B2(n1410), .ZN(n16) );
  AOI22_X1 U301 ( .A1(F[8]), .A2(n1428), .B1(E[8]), .B2(n1422), .ZN(n17) );
  NAND4_X1 U302 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U303 ( .A1(B[5]), .A2(n1403), .B1(A[5]), .B2(n1397), .ZN(n43) );
  AOI22_X1 U304 ( .A1(D[5]), .A2(n1415), .B1(C[5]), .B2(n1409), .ZN(n44) );
  AOI22_X1 U305 ( .A1(F[5]), .A2(n1427), .B1(E[5]), .B2(n1421), .ZN(n45) );
  NAND4_X1 U306 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U307 ( .A1(B[9]), .A2(n1404), .B1(A[9]), .B2(n1398), .ZN(n3) );
  AOI22_X1 U308 ( .A1(D[9]), .A2(n1416), .B1(C[9]), .B2(n1410), .ZN(n4) );
  AOI22_X1 U309 ( .A1(F[9]), .A2(n1428), .B1(E[9]), .B2(n1422), .ZN(n5) );
  NAND4_X1 U310 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U311 ( .A1(B[7]), .A2(n1404), .B1(A[7]), .B2(n1398), .ZN(n19) );
  AOI22_X1 U312 ( .A1(D[7]), .A2(n1416), .B1(C[7]), .B2(n1410), .ZN(n20) );
  AOI22_X1 U313 ( .A1(F[7]), .A2(n1428), .B1(E[7]), .B2(n1422), .ZN(n21) );
  NAND4_X1 U314 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U315 ( .A1(B[11]), .A2(n1399), .B1(A[11]), .B2(n1393), .ZN(n255) );
  AOI22_X1 U316 ( .A1(D[11]), .A2(n1411), .B1(C[11]), .B2(n1405), .ZN(n256) );
  AOI22_X1 U317 ( .A1(F[11]), .A2(n1423), .B1(E[11]), .B2(n1417), .ZN(n257) );
  NAND4_X1 U318 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U319 ( .A1(B[15]), .A2(n1399), .B1(A[15]), .B2(n1393), .ZN(n239) );
  AOI22_X1 U320 ( .A1(D[15]), .A2(n1411), .B1(C[15]), .B2(n1405), .ZN(n240) );
  AOI22_X1 U321 ( .A1(F[15]), .A2(n1423), .B1(E[15]), .B2(n1417), .ZN(n241) );
  NAND4_X1 U322 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U323 ( .A1(B[3]), .A2(n1401), .B1(A[3]), .B2(n1395), .ZN(n131) );
  AOI22_X1 U324 ( .A1(D[3]), .A2(n1413), .B1(C[3]), .B2(n1407), .ZN(n132) );
  AOI22_X1 U325 ( .A1(F[3]), .A2(n1425), .B1(E[3]), .B2(n1419), .ZN(n133) );
  NAND4_X1 U326 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U327 ( .A1(B[12]), .A2(n1399), .B1(A[12]), .B2(n1393), .ZN(n251) );
  AOI22_X1 U328 ( .A1(D[12]), .A2(n1411), .B1(C[12]), .B2(n1405), .ZN(n252) );
  AOI22_X1 U329 ( .A1(F[12]), .A2(n1423), .B1(E[12]), .B2(n1417), .ZN(n253) );
  NAND4_X1 U330 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U331 ( .A1(B[19]), .A2(n1399), .B1(A[19]), .B2(n1393), .ZN(n223) );
  AOI22_X1 U332 ( .A1(D[19]), .A2(n1411), .B1(C[19]), .B2(n1405), .ZN(n224) );
  AOI22_X1 U333 ( .A1(F[19]), .A2(n1423), .B1(E[19]), .B2(n1417), .ZN(n225) );
  NAND4_X1 U334 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U335 ( .A1(B[4]), .A2(n1402), .B1(A[4]), .B2(n1396), .ZN(n87) );
  AOI22_X1 U336 ( .A1(D[4]), .A2(n1414), .B1(C[4]), .B2(n1408), .ZN(n88) );
  AOI22_X1 U337 ( .A1(F[4]), .A2(n1426), .B1(E[4]), .B2(n1420), .ZN(n89) );
  NAND4_X1 U338 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U339 ( .A1(B[6]), .A2(n1404), .B1(A[6]), .B2(n1398), .ZN(n23) );
  AOI22_X1 U340 ( .A1(D[6]), .A2(n1416), .B1(C[6]), .B2(n1410), .ZN(n24) );
  AOI22_X1 U341 ( .A1(F[6]), .A2(n1428), .B1(E[6]), .B2(n1422), .ZN(n25) );
  NAND4_X1 U342 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U343 ( .A1(B[10]), .A2(n1399), .B1(A[10]), .B2(n1393), .ZN(n259) );
  AOI22_X1 U344 ( .A1(D[10]), .A2(n1411), .B1(C[10]), .B2(n1405), .ZN(n260) );
  AOI22_X1 U345 ( .A1(F[10]), .A2(n1423), .B1(E[10]), .B2(n1417), .ZN(n261) );
  NAND4_X1 U346 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U347 ( .A1(B[23]), .A2(n1400), .B1(A[23]), .B2(n1394), .ZN(n203) );
  AOI22_X1 U348 ( .A1(D[23]), .A2(n1412), .B1(C[23]), .B2(n1406), .ZN(n204) );
  AOI22_X1 U349 ( .A1(F[23]), .A2(n1424), .B1(E[23]), .B2(n1418), .ZN(n205) );
  NAND4_X1 U350 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U351 ( .A1(B[14]), .A2(n1399), .B1(A[14]), .B2(n1393), .ZN(n243) );
  AOI22_X1 U352 ( .A1(D[14]), .A2(n1411), .B1(C[14]), .B2(n1405), .ZN(n244) );
  AOI22_X1 U353 ( .A1(F[14]), .A2(n1423), .B1(E[14]), .B2(n1417), .ZN(n245) );
  NAND4_X1 U354 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U355 ( .A1(B[22]), .A2(n1400), .B1(A[22]), .B2(n1394), .ZN(n207) );
  AOI22_X1 U356 ( .A1(D[22]), .A2(n1412), .B1(C[22]), .B2(n1406), .ZN(n208) );
  AOI22_X1 U357 ( .A1(F[22]), .A2(n1424), .B1(E[22]), .B2(n1418), .ZN(n209) );
  NAND4_X1 U358 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U359 ( .A1(B[18]), .A2(n1399), .B1(A[18]), .B2(n1393), .ZN(n227) );
  AOI22_X1 U360 ( .A1(D[18]), .A2(n1411), .B1(C[18]), .B2(n1405), .ZN(n228) );
  AOI22_X1 U361 ( .A1(F[18]), .A2(n1423), .B1(E[18]), .B2(n1417), .ZN(n229) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1400), .B1(A[2]), .B2(n1394), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1412), .B1(C[2]), .B2(n1406), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1424), .B1(E[2]), .B2(n1418), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1399), .B1(A[1]), .B2(n1393), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1411), .B1(C[1]), .B2(n1405), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1423), .B1(E[1]), .B2(n1417), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1435), .B1(G[0]), .B2(n1429), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1398) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1404) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1410) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1416) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1422) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1428) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1434) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1440) );
endmodule


module MUX81_GENERIC_NBIT64_2 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444;

  BUF_X1 U1 ( .A(n13), .Z(n1402) );
  BUF_X1 U2 ( .A(n13), .Z(n1403) );
  BUF_X1 U3 ( .A(n12), .Z(n1408) );
  BUF_X1 U4 ( .A(n8), .Z(n1432) );
  BUF_X1 U5 ( .A(n8), .Z(n1433) );
  BUF_X1 U6 ( .A(n10), .Z(n1420) );
  BUF_X1 U7 ( .A(n10), .Z(n1421) );
  BUF_X1 U8 ( .A(n12), .Z(n1409) );
  BUF_X1 U9 ( .A(n13), .Z(n1404) );
  BUF_X1 U10 ( .A(n13), .Z(n1405) );
  BUF_X1 U11 ( .A(n12), .Z(n1410) );
  BUF_X1 U12 ( .A(n12), .Z(n1411) );
  BUF_X1 U13 ( .A(n10), .Z(n1422) );
  BUF_X1 U14 ( .A(n10), .Z(n1423) );
  BUF_X1 U15 ( .A(n8), .Z(n1434) );
  BUF_X1 U16 ( .A(n8), .Z(n1435) );
  BUF_X1 U17 ( .A(n11), .Z(n1416) );
  BUF_X1 U18 ( .A(n11), .Z(n1417) );
  BUF_X1 U19 ( .A(n11), .Z(n1414) );
  BUF_X1 U20 ( .A(n11), .Z(n1413) );
  BUF_X1 U21 ( .A(n13), .Z(n1401) );
  BUF_X1 U22 ( .A(n7), .Z(n1437) );
  BUF_X1 U23 ( .A(n7), .Z(n1438) );
  BUF_X1 U24 ( .A(n7), .Z(n1439) );
  BUF_X1 U25 ( .A(n9), .Z(n1428) );
  BUF_X1 U26 ( .A(n9), .Z(n1429) );
  BUF_X1 U27 ( .A(n7), .Z(n1440) );
  BUF_X1 U28 ( .A(n7), .Z(n1441) );
  BUF_X1 U29 ( .A(n9), .Z(n1426) );
  BUF_X1 U30 ( .A(n9), .Z(n1427) );
  BUF_X1 U31 ( .A(n9), .Z(n1425) );
  BUF_X1 U32 ( .A(n14), .Z(n1398) );
  BUF_X1 U33 ( .A(n14), .Z(n1399) );
  BUF_X1 U34 ( .A(n14), .Z(n1396) );
  BUF_X1 U35 ( .A(n14), .Z(n1397) );
  BUF_X1 U36 ( .A(n12), .Z(n1407) );
  BUF_X1 U37 ( .A(n14), .Z(n1395) );
  BUF_X1 U38 ( .A(n8), .Z(n1431) );
  BUF_X1 U39 ( .A(n10), .Z(n1419) );
  BUF_X1 U40 ( .A(n11), .Z(n1415) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1443), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1444), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1444), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1444), .A2(n1443), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1443) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1444) );
  NOR3_X1 U47 ( .A1(n1444), .A2(SEL[2]), .A3(n1443), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1443), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U52 ( .A1(B[59]), .A2(n1405), .B1(A[59]), .B2(n1399), .ZN(n47) );
  AOI22_X1 U53 ( .A1(D[59]), .A2(n1417), .B1(C[59]), .B2(n1411), .ZN(n48) );
  AOI22_X1 U54 ( .A1(H[59]), .A2(n1441), .B1(G[59]), .B2(n1435), .ZN(n50) );
  AOI22_X1 U55 ( .A1(F[59]), .A2(n1429), .B1(E[59]), .B2(n1423), .ZN(n49) );
  AOI22_X1 U56 ( .A1(F[41]), .A2(n1427), .B1(E[41]), .B2(n1421), .ZN(n125) );
  AOI22_X1 U57 ( .A1(F[62]), .A2(n1429), .B1(E[62]), .B2(n1423), .ZN(n33) );
  NAND4_X1 U58 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U59 ( .A1(B[49]), .A2(n1404), .B1(A[49]), .B2(n1398), .ZN(n91) );
  AOI22_X1 U60 ( .A1(D[49]), .A2(n1416), .B1(C[49]), .B2(n1410), .ZN(n92) );
  AOI22_X1 U61 ( .A1(H[49]), .A2(n1440), .B1(G[49]), .B2(n1434), .ZN(n94) );
  AOI22_X1 U62 ( .A1(F[51]), .A2(n1428), .B1(E[51]), .B2(n1422), .ZN(n81) );
  AOI22_X1 U63 ( .A1(F[37]), .A2(n1427), .B1(E[37]), .B2(n1421), .ZN(n145) );
  AOI22_X1 U64 ( .A1(F[33]), .A2(n1427), .B1(E[33]), .B2(n1421), .ZN(n161) );
  AOI22_X1 U65 ( .A1(F[57]), .A2(n1429), .B1(E[57]), .B2(n1423), .ZN(n57) );
  AOI22_X1 U66 ( .A1(F[61]), .A2(n1429), .B1(E[61]), .B2(n1423), .ZN(n37) );
  NAND4_X1 U67 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U68 ( .A1(B[52]), .A2(n1404), .B1(A[52]), .B2(n1398), .ZN(n75) );
  AOI22_X1 U69 ( .A1(D[52]), .A2(n1416), .B1(C[52]), .B2(n1410), .ZN(n76) );
  AOI22_X1 U70 ( .A1(H[52]), .A2(n1440), .B1(G[52]), .B2(n1434), .ZN(n78) );
  NAND4_X1 U71 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U72 ( .A1(B[38]), .A2(n1403), .B1(A[38]), .B2(n1397), .ZN(n139) );
  AOI22_X1 U73 ( .A1(D[38]), .A2(n1415), .B1(C[38]), .B2(n1409), .ZN(n140) );
  AOI22_X1 U74 ( .A1(H[38]), .A2(n1439), .B1(G[38]), .B2(n1433), .ZN(n142) );
  NAND4_X1 U75 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U76 ( .A1(H[29]), .A2(n1438), .B1(G[29]), .B2(n1432), .ZN(n182) );
  AOI22_X1 U77 ( .A1(B[29]), .A2(n1402), .B1(A[29]), .B2(n1396), .ZN(n179) );
  AOI22_X1 U78 ( .A1(D[29]), .A2(n1414), .B1(C[29]), .B2(n1408), .ZN(n180) );
  NAND4_X1 U79 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U80 ( .A1(B[46]), .A2(n1404), .B1(A[46]), .B2(n1398), .ZN(n103) );
  AOI22_X1 U81 ( .A1(D[46]), .A2(n1416), .B1(C[46]), .B2(n1410), .ZN(n104) );
  AOI22_X1 U82 ( .A1(H[46]), .A2(n1440), .B1(G[46]), .B2(n1434), .ZN(n106) );
  NAND4_X1 U83 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U84 ( .A1(B[53]), .A2(n1405), .B1(A[53]), .B2(n1399), .ZN(n71) );
  AOI22_X1 U85 ( .A1(D[53]), .A2(n1417), .B1(C[53]), .B2(n1411), .ZN(n72) );
  AOI22_X1 U86 ( .A1(H[53]), .A2(n1441), .B1(G[53]), .B2(n1435), .ZN(n74) );
  NAND4_X1 U87 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U88 ( .A1(B[56]), .A2(n1405), .B1(A[56]), .B2(n1399), .ZN(n59) );
  AOI22_X1 U89 ( .A1(D[56]), .A2(n1417), .B1(C[56]), .B2(n1411), .ZN(n60) );
  AOI22_X1 U90 ( .A1(H[56]), .A2(n1441), .B1(G[56]), .B2(n1435), .ZN(n62) );
  AOI22_X1 U91 ( .A1(F[29]), .A2(n1426), .B1(E[29]), .B2(n1420), .ZN(n181) );
  AOI22_X1 U92 ( .A1(F[28]), .A2(n1426), .B1(E[28]), .B2(n1420), .ZN(n185) );
  AOI22_X1 U93 ( .A1(F[39]), .A2(n1427), .B1(E[39]), .B2(n1421), .ZN(n137) );
  AOI22_X1 U94 ( .A1(F[38]), .A2(n1427), .B1(E[38]), .B2(n1421), .ZN(n141) );
  AOI22_X1 U95 ( .A1(F[43]), .A2(n1428), .B1(E[43]), .B2(n1422), .ZN(n117) );
  AOI22_X1 U96 ( .A1(F[31]), .A2(n1427), .B1(E[31]), .B2(n1421), .ZN(n169) );
  AOI22_X1 U97 ( .A1(F[40]), .A2(n1427), .B1(E[40]), .B2(n1421), .ZN(n129) );
  AOI22_X1 U98 ( .A1(F[35]), .A2(n1427), .B1(E[35]), .B2(n1421), .ZN(n153) );
  AOI22_X1 U99 ( .A1(F[44]), .A2(n1428), .B1(E[44]), .B2(n1422), .ZN(n113) );
  AOI22_X1 U100 ( .A1(F[32]), .A2(n1427), .B1(E[32]), .B2(n1421), .ZN(n165) );
  AOI22_X1 U101 ( .A1(F[45]), .A2(n1428), .B1(E[45]), .B2(n1422), .ZN(n109) );
  AOI22_X1 U102 ( .A1(F[47]), .A2(n1428), .B1(E[47]), .B2(n1422), .ZN(n101) );
  AOI22_X1 U103 ( .A1(F[48]), .A2(n1428), .B1(E[48]), .B2(n1422), .ZN(n97) );
  AOI22_X1 U104 ( .A1(F[49]), .A2(n1428), .B1(E[49]), .B2(n1422), .ZN(n93) );
  AOI22_X1 U105 ( .A1(F[55]), .A2(n1429), .B1(E[55]), .B2(n1423), .ZN(n65) );
  AOI22_X1 U106 ( .A1(F[30]), .A2(n1426), .B1(E[30]), .B2(n1420), .ZN(n173) );
  AOI22_X1 U107 ( .A1(F[53]), .A2(n1429), .B1(E[53]), .B2(n1423), .ZN(n73) );
  AOI22_X1 U108 ( .A1(F[56]), .A2(n1429), .B1(E[56]), .B2(n1423), .ZN(n61) );
  AOI22_X1 U109 ( .A1(F[54]), .A2(n1429), .B1(E[54]), .B2(n1423), .ZN(n69) );
  AOI22_X1 U110 ( .A1(F[34]), .A2(n1427), .B1(E[34]), .B2(n1421), .ZN(n157) );
  AOI22_X1 U111 ( .A1(F[63]), .A2(n1429), .B1(E[63]), .B2(n1423), .ZN(n29) );
  NAND4_X1 U112 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U113 ( .A1(B[50]), .A2(n1404), .B1(A[50]), .B2(n1398), .ZN(n83) );
  AOI22_X1 U114 ( .A1(D[50]), .A2(n1416), .B1(C[50]), .B2(n1410), .ZN(n84) );
  AOI22_X1 U115 ( .A1(H[50]), .A2(n1440), .B1(G[50]), .B2(n1434), .ZN(n86) );
  NAND4_X1 U116 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U117 ( .A1(B[57]), .A2(n1405), .B1(A[57]), .B2(n1399), .ZN(n55) );
  AOI22_X1 U118 ( .A1(D[57]), .A2(n1417), .B1(C[57]), .B2(n1411), .ZN(n56) );
  AOI22_X1 U119 ( .A1(H[57]), .A2(n1441), .B1(G[57]), .B2(n1435), .ZN(n58) );
  NAND4_X1 U120 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U121 ( .A1(B[47]), .A2(n1404), .B1(A[47]), .B2(n1398), .ZN(n99) );
  AOI22_X1 U122 ( .A1(D[47]), .A2(n1416), .B1(C[47]), .B2(n1410), .ZN(n100) );
  AOI22_X1 U123 ( .A1(H[47]), .A2(n1440), .B1(G[47]), .B2(n1434), .ZN(n102) );
  NAND4_X1 U124 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U125 ( .A1(B[54]), .A2(n1405), .B1(A[54]), .B2(n1399), .ZN(n67) );
  AOI22_X1 U126 ( .A1(D[54]), .A2(n1417), .B1(C[54]), .B2(n1411), .ZN(n68) );
  AOI22_X1 U127 ( .A1(H[54]), .A2(n1441), .B1(G[54]), .B2(n1435), .ZN(n70) );
  NAND4_X1 U128 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U129 ( .A1(B[48]), .A2(n1404), .B1(A[48]), .B2(n1398), .ZN(n95) );
  AOI22_X1 U130 ( .A1(D[48]), .A2(n1416), .B1(C[48]), .B2(n1410), .ZN(n96) );
  AOI22_X1 U131 ( .A1(H[48]), .A2(n1440), .B1(G[48]), .B2(n1434), .ZN(n98) );
  NAND4_X1 U132 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U133 ( .A1(B[58]), .A2(n1405), .B1(A[58]), .B2(n1399), .ZN(n51) );
  AOI22_X1 U134 ( .A1(D[58]), .A2(n1417), .B1(C[58]), .B2(n1411), .ZN(n52) );
  AOI22_X1 U135 ( .A1(H[58]), .A2(n1441), .B1(G[58]), .B2(n1435), .ZN(n54) );
  NAND4_X1 U136 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U137 ( .A1(H[32]), .A2(n1439), .B1(G[32]), .B2(n1433), .ZN(n166) );
  AOI22_X1 U138 ( .A1(B[32]), .A2(n1403), .B1(A[32]), .B2(n1397), .ZN(n163) );
  NAND4_X1 U139 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U140 ( .A1(B[61]), .A2(n1405), .B1(A[61]), .B2(n1399), .ZN(n35) );
  AOI22_X1 U141 ( .A1(D[61]), .A2(n1417), .B1(C[61]), .B2(n1411), .ZN(n36) );
  AOI22_X1 U142 ( .A1(H[61]), .A2(n1441), .B1(G[61]), .B2(n1435), .ZN(n38) );
  NAND4_X1 U143 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U144 ( .A1(D[28]), .A2(n1414), .B1(C[28]), .B2(n1408), .ZN(n184) );
  AOI22_X1 U145 ( .A1(H[28]), .A2(n1438), .B1(G[28]), .B2(n1432), .ZN(n186) );
  AOI22_X1 U146 ( .A1(B[28]), .A2(n1402), .B1(A[28]), .B2(n1396), .ZN(n183) );
  NAND4_X1 U147 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U148 ( .A1(B[37]), .A2(n1403), .B1(A[37]), .B2(n1397), .ZN(n143) );
  AOI22_X1 U149 ( .A1(D[37]), .A2(n1415), .B1(C[37]), .B2(n1409), .ZN(n144) );
  AOI22_X1 U150 ( .A1(H[37]), .A2(n1439), .B1(G[37]), .B2(n1433), .ZN(n146) );
  NAND4_X1 U151 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U152 ( .A1(B[36]), .A2(n1403), .B1(A[36]), .B2(n1397), .ZN(n147) );
  AOI22_X1 U153 ( .A1(D[36]), .A2(n1415), .B1(C[36]), .B2(n1409), .ZN(n148) );
  AOI22_X1 U154 ( .A1(H[36]), .A2(n1439), .B1(G[36]), .B2(n1433), .ZN(n150) );
  NAND4_X1 U155 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U156 ( .A1(B[41]), .A2(n1403), .B1(A[41]), .B2(n1397), .ZN(n123) );
  AOI22_X1 U157 ( .A1(D[41]), .A2(n1415), .B1(C[41]), .B2(n1409), .ZN(n124) );
  AOI22_X1 U158 ( .A1(H[41]), .A2(n1439), .B1(G[41]), .B2(n1433), .ZN(n126) );
  NAND4_X1 U159 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U160 ( .A1(B[40]), .A2(n1403), .B1(A[40]), .B2(n1397), .ZN(n127) );
  AOI22_X1 U161 ( .A1(D[40]), .A2(n1415), .B1(C[40]), .B2(n1409), .ZN(n128) );
  AOI22_X1 U162 ( .A1(H[40]), .A2(n1439), .B1(G[40]), .B2(n1433), .ZN(n130) );
  NAND4_X1 U163 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U164 ( .A1(B[44]), .A2(n1404), .B1(A[44]), .B2(n1398), .ZN(n111) );
  AOI22_X1 U165 ( .A1(D[44]), .A2(n1416), .B1(C[44]), .B2(n1410), .ZN(n112) );
  AOI22_X1 U166 ( .A1(H[44]), .A2(n1440), .B1(G[44]), .B2(n1434), .ZN(n114) );
  NAND4_X1 U167 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U168 ( .A1(B[33]), .A2(n1403), .B1(A[33]), .B2(n1397), .ZN(n159) );
  AOI22_X1 U169 ( .A1(H[33]), .A2(n1439), .B1(G[33]), .B2(n1433), .ZN(n162) );
  AOI22_X1 U170 ( .A1(D[33]), .A2(n1415), .B1(C[33]), .B2(n1409), .ZN(n160) );
  NAND4_X1 U171 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U172 ( .A1(B[45]), .A2(n1404), .B1(A[45]), .B2(n1398), .ZN(n107) );
  AOI22_X1 U173 ( .A1(D[45]), .A2(n1416), .B1(C[45]), .B2(n1410), .ZN(n108) );
  AOI22_X1 U174 ( .A1(H[45]), .A2(n1440), .B1(G[45]), .B2(n1434), .ZN(n110) );
  NAND4_X1 U175 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U176 ( .A1(H[30]), .A2(n1438), .B1(G[30]), .B2(n1432), .ZN(n174) );
  AOI22_X1 U177 ( .A1(B[30]), .A2(n1402), .B1(A[30]), .B2(n1396), .ZN(n171) );
  AOI22_X1 U178 ( .A1(D[30]), .A2(n1414), .B1(C[30]), .B2(n1408), .ZN(n172) );
  NAND4_X1 U179 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U180 ( .A1(H[31]), .A2(n1439), .B1(G[31]), .B2(n1433), .ZN(n170) );
  AOI22_X1 U181 ( .A1(B[31]), .A2(n1403), .B1(A[31]), .B2(n1397), .ZN(n167) );
  AOI22_X1 U182 ( .A1(D[31]), .A2(n1415), .B1(C[31]), .B2(n1409), .ZN(n168) );
  NAND4_X1 U183 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U184 ( .A1(B[35]), .A2(n1403), .B1(A[35]), .B2(n1397), .ZN(n151) );
  AOI22_X1 U185 ( .A1(D[35]), .A2(n1415), .B1(C[35]), .B2(n1409), .ZN(n152) );
  AOI22_X1 U186 ( .A1(H[35]), .A2(n1439), .B1(G[35]), .B2(n1433), .ZN(n154) );
  NAND4_X1 U187 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U188 ( .A1(B[34]), .A2(n1403), .B1(A[34]), .B2(n1397), .ZN(n155) );
  AOI22_X1 U189 ( .A1(H[34]), .A2(n1439), .B1(G[34]), .B2(n1433), .ZN(n158) );
  AOI22_X1 U190 ( .A1(D[34]), .A2(n1415), .B1(C[34]), .B2(n1409), .ZN(n156) );
  NAND4_X1 U191 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U192 ( .A1(B[42]), .A2(n1404), .B1(A[42]), .B2(n1398), .ZN(n119) );
  AOI22_X1 U193 ( .A1(D[42]), .A2(n1416), .B1(C[42]), .B2(n1410), .ZN(n120) );
  AOI22_X1 U194 ( .A1(H[42]), .A2(n1440), .B1(G[42]), .B2(n1434), .ZN(n122) );
  NAND4_X1 U195 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U196 ( .A1(B[60]), .A2(n1405), .B1(A[60]), .B2(n1399), .ZN(n39) );
  AOI22_X1 U197 ( .A1(D[60]), .A2(n1417), .B1(C[60]), .B2(n1411), .ZN(n40) );
  AOI22_X1 U198 ( .A1(H[60]), .A2(n1441), .B1(G[60]), .B2(n1435), .ZN(n42) );
  NAND4_X1 U199 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U200 ( .A1(B[51]), .A2(n1404), .B1(A[51]), .B2(n1398), .ZN(n79) );
  AOI22_X1 U201 ( .A1(D[51]), .A2(n1416), .B1(C[51]), .B2(n1410), .ZN(n80) );
  AOI22_X1 U202 ( .A1(H[51]), .A2(n1440), .B1(G[51]), .B2(n1434), .ZN(n82) );
  AOI22_X1 U203 ( .A1(F[60]), .A2(n1429), .B1(E[60]), .B2(n1423), .ZN(n41) );
  AOI22_X1 U204 ( .A1(F[52]), .A2(n1428), .B1(E[52]), .B2(n1422), .ZN(n77) );
  AOI22_X1 U205 ( .A1(F[36]), .A2(n1427), .B1(E[36]), .B2(n1421), .ZN(n149) );
  AOI22_X1 U206 ( .A1(F[42]), .A2(n1428), .B1(E[42]), .B2(n1422), .ZN(n121) );
  NAND4_X1 U207 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U208 ( .A1(B[39]), .A2(n1403), .B1(A[39]), .B2(n1397), .ZN(n135) );
  AOI22_X1 U209 ( .A1(D[39]), .A2(n1415), .B1(C[39]), .B2(n1409), .ZN(n136) );
  AOI22_X1 U210 ( .A1(H[39]), .A2(n1439), .B1(G[39]), .B2(n1433), .ZN(n138) );
  NAND4_X1 U211 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U212 ( .A1(B[55]), .A2(n1405), .B1(A[55]), .B2(n1399), .ZN(n63) );
  AOI22_X1 U213 ( .A1(D[55]), .A2(n1417), .B1(C[55]), .B2(n1411), .ZN(n64) );
  AOI22_X1 U214 ( .A1(H[55]), .A2(n1441), .B1(G[55]), .B2(n1435), .ZN(n66) );
  NAND4_X1 U215 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U216 ( .A1(B[43]), .A2(n1404), .B1(A[43]), .B2(n1398), .ZN(n115) );
  AOI22_X1 U217 ( .A1(D[43]), .A2(n1416), .B1(C[43]), .B2(n1410), .ZN(n116) );
  AOI22_X1 U218 ( .A1(H[43]), .A2(n1440), .B1(G[43]), .B2(n1434), .ZN(n118) );
  AOI22_X1 U219 ( .A1(F[46]), .A2(n1428), .B1(E[46]), .B2(n1422), .ZN(n105) );
  AOI22_X1 U220 ( .A1(F[50]), .A2(n1428), .B1(E[50]), .B2(n1422), .ZN(n85) );
  NAND4_X1 U221 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U222 ( .A1(B[62]), .A2(n1405), .B1(A[62]), .B2(n1399), .ZN(n31) );
  AOI22_X1 U223 ( .A1(D[62]), .A2(n1417), .B1(C[62]), .B2(n1411), .ZN(n32) );
  AOI22_X1 U224 ( .A1(H[62]), .A2(n1441), .B1(G[62]), .B2(n1435), .ZN(n34) );
  NAND4_X1 U225 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U226 ( .A1(B[63]), .A2(n1405), .B1(A[63]), .B2(n1399), .ZN(n27) );
  AOI22_X1 U227 ( .A1(D[63]), .A2(n1417), .B1(C[63]), .B2(n1411), .ZN(n28) );
  AOI22_X1 U228 ( .A1(H[63]), .A2(n1441), .B1(G[63]), .B2(n1435), .ZN(n30) );
  AOI22_X1 U229 ( .A1(F[58]), .A2(n1429), .B1(E[58]), .B2(n1423), .ZN(n53) );
  NAND4_X1 U230 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U231 ( .A1(B[0]), .A2(n1401), .B1(A[0]), .B2(n1395), .ZN(n263) );
  AOI22_X1 U232 ( .A1(D[0]), .A2(n1413), .B1(C[0]), .B2(n1407), .ZN(n264) );
  AOI22_X1 U233 ( .A1(F[0]), .A2(n1425), .B1(E[0]), .B2(n1419), .ZN(n265) );
  AOI22_X1 U234 ( .A1(H[13]), .A2(n1437), .B1(G[13]), .B2(n1431), .ZN(n250) );
  AOI22_X1 U235 ( .A1(H[17]), .A2(n1437), .B1(G[17]), .B2(n1431), .ZN(n234) );
  AOI22_X1 U236 ( .A1(H[21]), .A2(n1438), .B1(G[21]), .B2(n1432), .ZN(n214) );
  AOI22_X1 U237 ( .A1(H[25]), .A2(n1438), .B1(G[25]), .B2(n1432), .ZN(n198) );
  AOI22_X1 U238 ( .A1(H[5]), .A2(n1441), .B1(G[5]), .B2(n1435), .ZN(n46) );
  AOI22_X1 U239 ( .A1(H[9]), .A2(n1442), .B1(G[9]), .B2(n1436), .ZN(n6) );
  AOI22_X1 U240 ( .A1(H[7]), .A2(n1442), .B1(G[7]), .B2(n1436), .ZN(n22) );
  AOI22_X1 U241 ( .A1(H[11]), .A2(n1437), .B1(G[11]), .B2(n1431), .ZN(n258) );
  AOI22_X1 U242 ( .A1(H[15]), .A2(n1437), .B1(G[15]), .B2(n1431), .ZN(n242) );
  AOI22_X1 U243 ( .A1(H[23]), .A2(n1438), .B1(G[23]), .B2(n1432), .ZN(n206) );
  AOI22_X1 U244 ( .A1(H[27]), .A2(n1438), .B1(G[27]), .B2(n1432), .ZN(n190) );
  AOI22_X1 U245 ( .A1(H[19]), .A2(n1437), .B1(G[19]), .B2(n1431), .ZN(n226) );
  AOI22_X1 U246 ( .A1(H[3]), .A2(n1439), .B1(G[3]), .B2(n1433), .ZN(n134) );
  AOI22_X1 U247 ( .A1(H[20]), .A2(n1438), .B1(G[20]), .B2(n1432), .ZN(n218) );
  AOI22_X1 U248 ( .A1(H[12]), .A2(n1437), .B1(G[12]), .B2(n1431), .ZN(n254) );
  AOI22_X1 U249 ( .A1(H[4]), .A2(n1440), .B1(G[4]), .B2(n1434), .ZN(n90) );
  AOI22_X1 U250 ( .A1(H[8]), .A2(n1442), .B1(G[8]), .B2(n1436), .ZN(n18) );
  AOI22_X1 U251 ( .A1(H[24]), .A2(n1438), .B1(G[24]), .B2(n1432), .ZN(n202) );
  AOI22_X1 U252 ( .A1(H[16]), .A2(n1437), .B1(G[16]), .B2(n1431), .ZN(n238) );
  AOI22_X1 U253 ( .A1(H[6]), .A2(n1442), .B1(G[6]), .B2(n1436), .ZN(n26) );
  AOI22_X1 U254 ( .A1(H[10]), .A2(n1437), .B1(G[10]), .B2(n1431), .ZN(n262) );
  AOI22_X1 U255 ( .A1(H[14]), .A2(n1437), .B1(G[14]), .B2(n1431), .ZN(n246) );
  AOI22_X1 U256 ( .A1(H[22]), .A2(n1438), .B1(G[22]), .B2(n1432), .ZN(n210) );
  AOI22_X1 U257 ( .A1(H[26]), .A2(n1438), .B1(G[26]), .B2(n1432), .ZN(n194) );
  AOI22_X1 U258 ( .A1(H[18]), .A2(n1437), .B1(G[18]), .B2(n1431), .ZN(n230) );
  AOI22_X1 U259 ( .A1(H[2]), .A2(n1438), .B1(G[2]), .B2(n1432), .ZN(n178) );
  AOI22_X1 U260 ( .A1(H[1]), .A2(n1437), .B1(G[1]), .B2(n1431), .ZN(n222) );
  NAND4_X1 U261 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U262 ( .A1(B[13]), .A2(n1401), .B1(A[13]), .B2(n1395), .ZN(n247) );
  AOI22_X1 U263 ( .A1(D[13]), .A2(n1413), .B1(C[13]), .B2(n1407), .ZN(n248) );
  AOI22_X1 U264 ( .A1(F[13]), .A2(n1425), .B1(E[13]), .B2(n1419), .ZN(n249) );
  NAND4_X1 U265 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U266 ( .A1(B[17]), .A2(n1401), .B1(A[17]), .B2(n1395), .ZN(n231) );
  AOI22_X1 U267 ( .A1(D[17]), .A2(n1413), .B1(C[17]), .B2(n1407), .ZN(n232) );
  AOI22_X1 U268 ( .A1(F[17]), .A2(n1425), .B1(E[17]), .B2(n1419), .ZN(n233) );
  NAND4_X1 U269 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U270 ( .A1(B[12]), .A2(n1401), .B1(A[12]), .B2(n1395), .ZN(n251) );
  AOI22_X1 U271 ( .A1(D[12]), .A2(n1413), .B1(C[12]), .B2(n1407), .ZN(n252) );
  AOI22_X1 U272 ( .A1(F[12]), .A2(n1425), .B1(E[12]), .B2(n1419), .ZN(n253) );
  NAND4_X1 U273 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U274 ( .A1(B[21]), .A2(n1402), .B1(A[21]), .B2(n1396), .ZN(n211) );
  AOI22_X1 U275 ( .A1(D[21]), .A2(n1414), .B1(C[21]), .B2(n1408), .ZN(n212) );
  AOI22_X1 U276 ( .A1(F[21]), .A2(n1426), .B1(E[21]), .B2(n1420), .ZN(n213) );
  NAND4_X1 U277 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U278 ( .A1(B[5]), .A2(n1405), .B1(A[5]), .B2(n1399), .ZN(n43) );
  AOI22_X1 U279 ( .A1(D[5]), .A2(n1417), .B1(C[5]), .B2(n1411), .ZN(n44) );
  AOI22_X1 U280 ( .A1(F[5]), .A2(n1429), .B1(E[5]), .B2(n1423), .ZN(n45) );
  NAND4_X1 U281 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U282 ( .A1(B[7]), .A2(n1406), .B1(A[7]), .B2(n1400), .ZN(n19) );
  AOI22_X1 U283 ( .A1(D[7]), .A2(n1418), .B1(C[7]), .B2(n1412), .ZN(n20) );
  AOI22_X1 U284 ( .A1(F[7]), .A2(n1430), .B1(E[7]), .B2(n1424), .ZN(n21) );
  NAND4_X1 U285 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U286 ( .A1(B[11]), .A2(n1401), .B1(A[11]), .B2(n1395), .ZN(n255) );
  AOI22_X1 U287 ( .A1(D[11]), .A2(n1413), .B1(C[11]), .B2(n1407), .ZN(n256) );
  AOI22_X1 U288 ( .A1(F[11]), .A2(n1425), .B1(E[11]), .B2(n1419), .ZN(n257) );
  NAND4_X1 U289 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U290 ( .A1(B[23]), .A2(n1402), .B1(A[23]), .B2(n1396), .ZN(n203) );
  AOI22_X1 U291 ( .A1(D[23]), .A2(n1414), .B1(C[23]), .B2(n1408), .ZN(n204) );
  AOI22_X1 U292 ( .A1(F[23]), .A2(n1426), .B1(E[23]), .B2(n1420), .ZN(n205) );
  NAND4_X1 U293 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U294 ( .A1(B[27]), .A2(n1402), .B1(A[27]), .B2(n1396), .ZN(n187) );
  AOI22_X1 U295 ( .A1(D[27]), .A2(n1414), .B1(C[27]), .B2(n1408), .ZN(n188) );
  AOI22_X1 U296 ( .A1(F[27]), .A2(n1426), .B1(E[27]), .B2(n1420), .ZN(n189) );
  NAND4_X1 U297 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U298 ( .A1(B[3]), .A2(n1403), .B1(A[3]), .B2(n1397), .ZN(n131) );
  AOI22_X1 U299 ( .A1(D[3]), .A2(n1415), .B1(C[3]), .B2(n1409), .ZN(n132) );
  AOI22_X1 U300 ( .A1(F[3]), .A2(n1427), .B1(E[3]), .B2(n1421), .ZN(n133) );
  NAND4_X1 U301 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U302 ( .A1(B[20]), .A2(n1402), .B1(A[20]), .B2(n1396), .ZN(n215) );
  AOI22_X1 U303 ( .A1(D[20]), .A2(n1414), .B1(C[20]), .B2(n1408), .ZN(n216) );
  AOI22_X1 U304 ( .A1(F[20]), .A2(n1426), .B1(E[20]), .B2(n1420), .ZN(n217) );
  NAND4_X1 U305 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U306 ( .A1(B[25]), .A2(n1402), .B1(A[25]), .B2(n1396), .ZN(n195) );
  AOI22_X1 U307 ( .A1(D[25]), .A2(n1414), .B1(C[25]), .B2(n1408), .ZN(n196) );
  AOI22_X1 U308 ( .A1(F[25]), .A2(n1426), .B1(E[25]), .B2(n1420), .ZN(n197) );
  NAND4_X1 U309 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U310 ( .A1(B[9]), .A2(n1406), .B1(A[9]), .B2(n1400), .ZN(n3) );
  AOI22_X1 U311 ( .A1(D[9]), .A2(n1418), .B1(C[9]), .B2(n1412), .ZN(n4) );
  AOI22_X1 U312 ( .A1(F[9]), .A2(n1430), .B1(E[9]), .B2(n1424), .ZN(n5) );
  NAND4_X1 U313 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U314 ( .A1(B[8]), .A2(n1406), .B1(A[8]), .B2(n1400), .ZN(n15) );
  AOI22_X1 U315 ( .A1(D[8]), .A2(n1418), .B1(C[8]), .B2(n1412), .ZN(n16) );
  AOI22_X1 U316 ( .A1(F[8]), .A2(n1430), .B1(E[8]), .B2(n1424), .ZN(n17) );
  NAND4_X1 U317 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U318 ( .A1(B[4]), .A2(n1404), .B1(A[4]), .B2(n1398), .ZN(n87) );
  AOI22_X1 U319 ( .A1(D[4]), .A2(n1416), .B1(C[4]), .B2(n1410), .ZN(n88) );
  AOI22_X1 U320 ( .A1(F[4]), .A2(n1428), .B1(E[4]), .B2(n1422), .ZN(n89) );
  NAND4_X1 U321 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U322 ( .A1(B[24]), .A2(n1402), .B1(A[24]), .B2(n1396), .ZN(n199) );
  AOI22_X1 U323 ( .A1(D[24]), .A2(n1414), .B1(C[24]), .B2(n1408), .ZN(n200) );
  AOI22_X1 U324 ( .A1(F[24]), .A2(n1426), .B1(E[24]), .B2(n1420), .ZN(n201) );
  NAND4_X1 U325 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U326 ( .A1(B[15]), .A2(n1401), .B1(A[15]), .B2(n1395), .ZN(n239) );
  AOI22_X1 U327 ( .A1(D[15]), .A2(n1413), .B1(C[15]), .B2(n1407), .ZN(n240) );
  AOI22_X1 U328 ( .A1(F[15]), .A2(n1425), .B1(E[15]), .B2(n1419), .ZN(n241) );
  NAND4_X1 U329 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U330 ( .A1(B[19]), .A2(n1401), .B1(A[19]), .B2(n1395), .ZN(n223) );
  AOI22_X1 U331 ( .A1(D[19]), .A2(n1413), .B1(C[19]), .B2(n1407), .ZN(n224) );
  AOI22_X1 U332 ( .A1(F[19]), .A2(n1425), .B1(E[19]), .B2(n1419), .ZN(n225) );
  NAND4_X1 U333 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U334 ( .A1(B[6]), .A2(n1406), .B1(A[6]), .B2(n1400), .ZN(n23) );
  AOI22_X1 U335 ( .A1(D[6]), .A2(n1418), .B1(C[6]), .B2(n1412), .ZN(n24) );
  AOI22_X1 U336 ( .A1(F[6]), .A2(n1430), .B1(E[6]), .B2(n1424), .ZN(n25) );
  NAND4_X1 U337 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U338 ( .A1(B[10]), .A2(n1401), .B1(A[10]), .B2(n1395), .ZN(n259) );
  AOI22_X1 U339 ( .A1(D[10]), .A2(n1413), .B1(C[10]), .B2(n1407), .ZN(n260) );
  AOI22_X1 U340 ( .A1(F[10]), .A2(n1425), .B1(E[10]), .B2(n1419), .ZN(n261) );
  NAND4_X1 U341 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U342 ( .A1(B[16]), .A2(n1401), .B1(A[16]), .B2(n1395), .ZN(n235) );
  AOI22_X1 U343 ( .A1(D[16]), .A2(n1413), .B1(C[16]), .B2(n1407), .ZN(n236) );
  AOI22_X1 U344 ( .A1(F[16]), .A2(n1425), .B1(E[16]), .B2(n1419), .ZN(n237) );
  NAND4_X1 U345 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U346 ( .A1(B[14]), .A2(n1401), .B1(A[14]), .B2(n1395), .ZN(n243) );
  AOI22_X1 U347 ( .A1(D[14]), .A2(n1413), .B1(C[14]), .B2(n1407), .ZN(n244) );
  AOI22_X1 U348 ( .A1(F[14]), .A2(n1425), .B1(E[14]), .B2(n1419), .ZN(n245) );
  NAND4_X1 U349 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U350 ( .A1(B[22]), .A2(n1402), .B1(A[22]), .B2(n1396), .ZN(n207) );
  AOI22_X1 U351 ( .A1(D[22]), .A2(n1414), .B1(C[22]), .B2(n1408), .ZN(n208) );
  AOI22_X1 U352 ( .A1(F[22]), .A2(n1426), .B1(E[22]), .B2(n1420), .ZN(n209) );
  NAND4_X1 U353 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U354 ( .A1(B[26]), .A2(n1402), .B1(A[26]), .B2(n1396), .ZN(n191) );
  AOI22_X1 U355 ( .A1(D[26]), .A2(n1414), .B1(C[26]), .B2(n1408), .ZN(n192) );
  AOI22_X1 U356 ( .A1(F[26]), .A2(n1426), .B1(E[26]), .B2(n1420), .ZN(n193) );
  NAND4_X1 U357 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U358 ( .A1(B[18]), .A2(n1401), .B1(A[18]), .B2(n1395), .ZN(n227) );
  AOI22_X1 U359 ( .A1(D[18]), .A2(n1413), .B1(C[18]), .B2(n1407), .ZN(n228) );
  AOI22_X1 U360 ( .A1(F[18]), .A2(n1425), .B1(E[18]), .B2(n1419), .ZN(n229) );
  NAND4_X1 U361 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U362 ( .A1(B[2]), .A2(n1402), .B1(A[2]), .B2(n1396), .ZN(n175) );
  AOI22_X1 U363 ( .A1(D[2]), .A2(n1414), .B1(C[2]), .B2(n1408), .ZN(n176) );
  AOI22_X1 U364 ( .A1(F[2]), .A2(n1426), .B1(E[2]), .B2(n1420), .ZN(n177) );
  NAND4_X1 U365 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U366 ( .A1(B[1]), .A2(n1401), .B1(A[1]), .B2(n1395), .ZN(n219) );
  AOI22_X1 U367 ( .A1(D[1]), .A2(n1413), .B1(C[1]), .B2(n1407), .ZN(n220) );
  AOI22_X1 U368 ( .A1(F[1]), .A2(n1425), .B1(E[1]), .B2(n1419), .ZN(n221) );
  AOI22_X1 U369 ( .A1(H[0]), .A2(n1437), .B1(G[0]), .B2(n1431), .ZN(n266) );
  AOI22_X1 U370 ( .A1(D[32]), .A2(n1415), .B1(C[32]), .B2(n1409), .ZN(n164) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1400) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1406) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1412) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1418) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1424) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1430) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1436) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1442) );
endmodule


module MUX81_GENERIC_NBIT64_1 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [63:0] F;
  input [63:0] G;
  input [63:0] H;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444;

  BUF_X1 U1 ( .A(n13), .Z(n1404) );
  BUF_X1 U2 ( .A(n13), .Z(n1405) );
  BUF_X1 U3 ( .A(n13), .Z(n1402) );
  BUF_X1 U4 ( .A(n13), .Z(n1403) );
  BUF_X1 U5 ( .A(n12), .Z(n1410) );
  BUF_X1 U6 ( .A(n12), .Z(n1411) );
  BUF_X1 U7 ( .A(n12), .Z(n1409) );
  BUF_X1 U8 ( .A(n10), .Z(n1422) );
  BUF_X1 U9 ( .A(n8), .Z(n1434) );
  BUF_X1 U10 ( .A(n10), .Z(n1423) );
  BUF_X1 U11 ( .A(n8), .Z(n1435) );
  BUF_X1 U12 ( .A(n8), .Z(n1433) );
  BUF_X1 U13 ( .A(n10), .Z(n1420) );
  BUF_X1 U14 ( .A(n10), .Z(n1421) );
  BUF_X1 U15 ( .A(n11), .Z(n1416) );
  BUF_X1 U16 ( .A(n11), .Z(n1417) );
  BUF_X1 U17 ( .A(n11), .Z(n1414) );
  BUF_X1 U18 ( .A(n11), .Z(n1415) );
  BUF_X1 U19 ( .A(n11), .Z(n1413) );
  BUF_X1 U20 ( .A(n13), .Z(n1401) );
  BUF_X1 U21 ( .A(n7), .Z(n1437) );
  BUF_X1 U22 ( .A(n7), .Z(n1438) );
  BUF_X1 U23 ( .A(n9), .Z(n1428) );
  BUF_X1 U24 ( .A(n7), .Z(n1440) );
  BUF_X1 U25 ( .A(n9), .Z(n1429) );
  BUF_X1 U26 ( .A(n7), .Z(n1441) );
  BUF_X1 U27 ( .A(n7), .Z(n1439) );
  BUF_X1 U28 ( .A(n9), .Z(n1426) );
  BUF_X1 U29 ( .A(n9), .Z(n1427) );
  BUF_X1 U30 ( .A(n9), .Z(n1425) );
  BUF_X1 U31 ( .A(n14), .Z(n1398) );
  BUF_X1 U32 ( .A(n14), .Z(n1399) );
  BUF_X1 U33 ( .A(n12), .Z(n1408) );
  BUF_X1 U34 ( .A(n14), .Z(n1396) );
  BUF_X1 U35 ( .A(n14), .Z(n1397) );
  BUF_X1 U36 ( .A(n12), .Z(n1407) );
  BUF_X1 U37 ( .A(n14), .Z(n1395) );
  BUF_X1 U38 ( .A(n8), .Z(n1431) );
  BUF_X1 U39 ( .A(n8), .Z(n1432) );
  BUF_X1 U40 ( .A(n10), .Z(n1419) );
  NOR3_X1 U41 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n1443), .ZN(n12) );
  NOR3_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n1444), .ZN(n13) );
  AND3_X1 U43 ( .A1(SEL[1]), .A2(n1444), .A3(SEL[2]), .ZN(n8) );
  AND3_X1 U44 ( .A1(n1444), .A2(n1443), .A3(SEL[2]), .ZN(n10) );
  INV_X1 U45 ( .A(SEL[1]), .ZN(n1443) );
  INV_X1 U46 ( .A(SEL[0]), .ZN(n1444) );
  NOR3_X1 U47 ( .A1(n1444), .A2(SEL[2]), .A3(n1443), .ZN(n11) );
  NOR3_X1 U48 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n14) );
  AND3_X1 U49 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n7) );
  AND3_X1 U50 ( .A1(SEL[0]), .A2(n1443), .A3(SEL[2]), .ZN(n9) );
  NAND4_X1 U51 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[54]) );
  AOI22_X1 U52 ( .A1(B[54]), .A2(n1405), .B1(A[54]), .B2(n1399), .ZN(n67) );
  AOI22_X1 U53 ( .A1(D[54]), .A2(n1417), .B1(C[54]), .B2(n1411), .ZN(n68) );
  AOI22_X1 U54 ( .A1(H[54]), .A2(n1441), .B1(G[54]), .B2(n1435), .ZN(n70) );
  AOI22_X1 U55 ( .A1(F[62]), .A2(n1429), .B1(E[62]), .B2(n1423), .ZN(n33) );
  AOI22_X1 U56 ( .A1(F[59]), .A2(n1429), .B1(E[59]), .B2(n1423), .ZN(n49) );
  NAND4_X1 U57 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(Y[58]) );
  AOI22_X1 U58 ( .A1(B[58]), .A2(n1405), .B1(A[58]), .B2(n1399), .ZN(n51) );
  AOI22_X1 U59 ( .A1(D[58]), .A2(n1417), .B1(C[58]), .B2(n1411), .ZN(n52) );
  AOI22_X1 U60 ( .A1(H[58]), .A2(n1441), .B1(G[58]), .B2(n1435), .ZN(n54) );
  NAND4_X1 U61 ( .A1(n59), .A2(n60), .A3(n61), .A4(n62), .ZN(Y[56]) );
  AOI22_X1 U62 ( .A1(B[56]), .A2(n1405), .B1(A[56]), .B2(n1399), .ZN(n59) );
  AOI22_X1 U63 ( .A1(D[56]), .A2(n1417), .B1(C[56]), .B2(n1411), .ZN(n60) );
  AOI22_X1 U64 ( .A1(H[56]), .A2(n1441), .B1(G[56]), .B2(n1435), .ZN(n62) );
  NAND4_X1 U65 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .ZN(Y[50]) );
  AOI22_X1 U66 ( .A1(B[50]), .A2(n1404), .B1(A[50]), .B2(n1398), .ZN(n83) );
  AOI22_X1 U67 ( .A1(D[50]), .A2(n1416), .B1(C[50]), .B2(n1410), .ZN(n84) );
  AOI22_X1 U68 ( .A1(H[50]), .A2(n1440), .B1(G[50]), .B2(n1434), .ZN(n86) );
  NAND4_X1 U69 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .ZN(Y[47]) );
  AOI22_X1 U70 ( .A1(B[47]), .A2(n1404), .B1(A[47]), .B2(n1398), .ZN(n99) );
  AOI22_X1 U71 ( .A1(D[47]), .A2(n1416), .B1(C[47]), .B2(n1410), .ZN(n100) );
  AOI22_X1 U72 ( .A1(H[47]), .A2(n1440), .B1(G[47]), .B2(n1434), .ZN(n102) );
  NAND4_X1 U73 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(Y[57]) );
  AOI22_X1 U74 ( .A1(B[57]), .A2(n1405), .B1(A[57]), .B2(n1399), .ZN(n55) );
  AOI22_X1 U75 ( .A1(D[57]), .A2(n1417), .B1(C[57]), .B2(n1411), .ZN(n56) );
  AOI22_X1 U76 ( .A1(H[57]), .A2(n1441), .B1(G[57]), .B2(n1435), .ZN(n58) );
  AOI22_X1 U77 ( .A1(F[47]), .A2(n1428), .B1(E[47]), .B2(n1422), .ZN(n101) );
  AOI22_X1 U78 ( .A1(F[51]), .A2(n1428), .B1(E[51]), .B2(n1422), .ZN(n81) );
  AOI22_X1 U79 ( .A1(F[55]), .A2(n1429), .B1(E[55]), .B2(n1423), .ZN(n65) );
  AOI22_X1 U80 ( .A1(F[57]), .A2(n1429), .B1(E[57]), .B2(n1423), .ZN(n57) );
  AOI22_X1 U81 ( .A1(F[49]), .A2(n1428), .B1(E[49]), .B2(n1422), .ZN(n93) );
  AOI22_X1 U82 ( .A1(F[52]), .A2(n1428), .B1(E[52]), .B2(n1422), .ZN(n77) );
  AOI22_X1 U83 ( .A1(F[41]), .A2(n1427), .B1(E[41]), .B2(n1421), .ZN(n125) );
  AOI22_X1 U84 ( .A1(F[42]), .A2(n1428), .B1(E[42]), .B2(n1422), .ZN(n121) );
  AOI22_X1 U85 ( .A1(F[43]), .A2(n1428), .B1(E[43]), .B2(n1422), .ZN(n117) );
  AOI22_X1 U86 ( .A1(F[45]), .A2(n1428), .B1(E[45]), .B2(n1422), .ZN(n109) );
  AOI22_X1 U87 ( .A1(F[53]), .A2(n1429), .B1(E[53]), .B2(n1423), .ZN(n73) );
  AOI22_X1 U88 ( .A1(F[63]), .A2(n1429), .B1(E[63]), .B2(n1423), .ZN(n29) );
  NAND4_X1 U89 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(Y[62]) );
  AOI22_X1 U90 ( .A1(B[62]), .A2(n1405), .B1(A[62]), .B2(n1399), .ZN(n31) );
  AOI22_X1 U91 ( .A1(D[62]), .A2(n1417), .B1(C[62]), .B2(n1411), .ZN(n32) );
  AOI22_X1 U92 ( .A1(H[62]), .A2(n1441), .B1(G[62]), .B2(n1435), .ZN(n34) );
  NAND4_X1 U93 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(Y[60]) );
  AOI22_X1 U94 ( .A1(B[60]), .A2(n1405), .B1(A[60]), .B2(n1399), .ZN(n39) );
  AOI22_X1 U95 ( .A1(D[60]), .A2(n1417), .B1(C[60]), .B2(n1411), .ZN(n40) );
  AOI22_X1 U96 ( .A1(H[60]), .A2(n1441), .B1(G[60]), .B2(n1435), .ZN(n42) );
  NAND4_X1 U97 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(Y[61]) );
  AOI22_X1 U98 ( .A1(B[61]), .A2(n1405), .B1(A[61]), .B2(n1399), .ZN(n35) );
  AOI22_X1 U99 ( .A1(D[61]), .A2(n1417), .B1(C[61]), .B2(n1411), .ZN(n36) );
  AOI22_X1 U100 ( .A1(H[61]), .A2(n1441), .B1(G[61]), .B2(n1435), .ZN(n38) );
  NAND4_X1 U101 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(Y[48]) );
  AOI22_X1 U102 ( .A1(B[48]), .A2(n1404), .B1(A[48]), .B2(n1398), .ZN(n95) );
  AOI22_X1 U103 ( .A1(D[48]), .A2(n1416), .B1(C[48]), .B2(n1410), .ZN(n96) );
  AOI22_X1 U104 ( .A1(H[48]), .A2(n1440), .B1(G[48]), .B2(n1434), .ZN(n98) );
  NAND4_X1 U105 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(Y[49]) );
  AOI22_X1 U106 ( .A1(B[49]), .A2(n1404), .B1(A[49]), .B2(n1398), .ZN(n91) );
  AOI22_X1 U107 ( .A1(D[49]), .A2(n1416), .B1(C[49]), .B2(n1410), .ZN(n92) );
  AOI22_X1 U108 ( .A1(H[49]), .A2(n1440), .B1(G[49]), .B2(n1434), .ZN(n94) );
  NAND4_X1 U109 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(Y[52]) );
  AOI22_X1 U110 ( .A1(B[52]), .A2(n1404), .B1(A[52]), .B2(n1398), .ZN(n75) );
  AOI22_X1 U111 ( .A1(D[52]), .A2(n1416), .B1(C[52]), .B2(n1410), .ZN(n76) );
  AOI22_X1 U112 ( .A1(H[52]), .A2(n1440), .B1(G[52]), .B2(n1434), .ZN(n78) );
  NAND4_X1 U113 ( .A1(n123), .A2(n124), .A3(n125), .A4(n126), .ZN(Y[41]) );
  AOI22_X1 U114 ( .A1(B[41]), .A2(n1403), .B1(A[41]), .B2(n1397), .ZN(n123) );
  AOI22_X1 U115 ( .A1(D[41]), .A2(n1415), .B1(C[41]), .B2(n1409), .ZN(n124) );
  AOI22_X1 U116 ( .A1(H[41]), .A2(n1439), .B1(G[41]), .B2(n1433), .ZN(n126) );
  NAND4_X1 U117 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(Y[42]) );
  AOI22_X1 U118 ( .A1(B[42]), .A2(n1404), .B1(A[42]), .B2(n1398), .ZN(n119) );
  AOI22_X1 U119 ( .A1(D[42]), .A2(n1416), .B1(C[42]), .B2(n1410), .ZN(n120) );
  AOI22_X1 U120 ( .A1(H[42]), .A2(n1440), .B1(G[42]), .B2(n1434), .ZN(n122) );
  NAND4_X1 U121 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(Y[44]) );
  AOI22_X1 U122 ( .A1(B[44]), .A2(n1404), .B1(A[44]), .B2(n1398), .ZN(n111) );
  AOI22_X1 U123 ( .A1(D[44]), .A2(n1416), .B1(C[44]), .B2(n1410), .ZN(n112) );
  AOI22_X1 U124 ( .A1(H[44]), .A2(n1440), .B1(G[44]), .B2(n1434), .ZN(n114) );
  NAND4_X1 U125 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(Y[45]) );
  AOI22_X1 U126 ( .A1(B[45]), .A2(n1404), .B1(A[45]), .B2(n1398), .ZN(n107) );
  AOI22_X1 U127 ( .A1(D[45]), .A2(n1416), .B1(C[45]), .B2(n1410), .ZN(n108) );
  AOI22_X1 U128 ( .A1(H[45]), .A2(n1440), .B1(G[45]), .B2(n1434), .ZN(n110) );
  NAND4_X1 U129 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(Y[51]) );
  AOI22_X1 U130 ( .A1(B[51]), .A2(n1404), .B1(A[51]), .B2(n1398), .ZN(n79) );
  AOI22_X1 U131 ( .A1(D[51]), .A2(n1416), .B1(C[51]), .B2(n1410), .ZN(n80) );
  AOI22_X1 U132 ( .A1(H[51]), .A2(n1440), .B1(G[51]), .B2(n1434), .ZN(n82) );
  NAND4_X1 U133 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(Y[46]) );
  AOI22_X1 U134 ( .A1(B[46]), .A2(n1404), .B1(A[46]), .B2(n1398), .ZN(n103) );
  AOI22_X1 U135 ( .A1(D[46]), .A2(n1416), .B1(C[46]), .B2(n1410), .ZN(n104) );
  AOI22_X1 U136 ( .A1(H[46]), .A2(n1440), .B1(G[46]), .B2(n1434), .ZN(n106) );
  NAND4_X1 U137 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(Y[53]) );
  AOI22_X1 U138 ( .A1(B[53]), .A2(n1405), .B1(A[53]), .B2(n1399), .ZN(n71) );
  AOI22_X1 U139 ( .A1(D[53]), .A2(n1417), .B1(C[53]), .B2(n1411), .ZN(n72) );
  AOI22_X1 U140 ( .A1(H[53]), .A2(n1441), .B1(G[53]), .B2(n1435), .ZN(n74) );
  NAND4_X1 U141 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(Y[55]) );
  AOI22_X1 U142 ( .A1(B[55]), .A2(n1405), .B1(A[55]), .B2(n1399), .ZN(n63) );
  AOI22_X1 U143 ( .A1(D[55]), .A2(n1417), .B1(C[55]), .B2(n1411), .ZN(n64) );
  AOI22_X1 U144 ( .A1(H[55]), .A2(n1441), .B1(G[55]), .B2(n1435), .ZN(n66) );
  AOI22_X1 U145 ( .A1(F[48]), .A2(n1428), .B1(E[48]), .B2(n1422), .ZN(n97) );
  AOI22_X1 U146 ( .A1(F[44]), .A2(n1428), .B1(E[44]), .B2(n1422), .ZN(n113) );
  AOI22_X1 U147 ( .A1(F[60]), .A2(n1429), .B1(E[60]), .B2(n1423), .ZN(n41) );
  AOI22_X1 U148 ( .A1(F[56]), .A2(n1429), .B1(E[56]), .B2(n1423), .ZN(n61) );
  AOI22_X1 U149 ( .A1(F[50]), .A2(n1428), .B1(E[50]), .B2(n1422), .ZN(n85) );
  AOI22_X1 U150 ( .A1(F[46]), .A2(n1428), .B1(E[46]), .B2(n1422), .ZN(n105) );
  NAND4_X1 U151 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(Y[43]) );
  AOI22_X1 U152 ( .A1(B[43]), .A2(n1404), .B1(A[43]), .B2(n1398), .ZN(n115) );
  AOI22_X1 U153 ( .A1(D[43]), .A2(n1416), .B1(C[43]), .B2(n1410), .ZN(n116) );
  AOI22_X1 U154 ( .A1(H[43]), .A2(n1440), .B1(G[43]), .B2(n1434), .ZN(n118) );
  NAND4_X1 U155 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(Y[59]) );
  AOI22_X1 U156 ( .A1(B[59]), .A2(n1405), .B1(A[59]), .B2(n1399), .ZN(n47) );
  AOI22_X1 U157 ( .A1(D[59]), .A2(n1417), .B1(C[59]), .B2(n1411), .ZN(n48) );
  AOI22_X1 U158 ( .A1(H[59]), .A2(n1441), .B1(G[59]), .B2(n1435), .ZN(n50) );
  AOI22_X1 U159 ( .A1(F[54]), .A2(n1429), .B1(E[54]), .B2(n1423), .ZN(n69) );
  AOI22_X1 U160 ( .A1(F[61]), .A2(n1429), .B1(E[61]), .B2(n1423), .ZN(n37) );
  AOI22_X1 U161 ( .A1(F[58]), .A2(n1429), .B1(E[58]), .B2(n1423), .ZN(n53) );
  NAND4_X1 U162 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(Y[63]) );
  AOI22_X1 U163 ( .A1(B[63]), .A2(n1405), .B1(A[63]), .B2(n1399), .ZN(n27) );
  AOI22_X1 U164 ( .A1(D[63]), .A2(n1417), .B1(C[63]), .B2(n1411), .ZN(n28) );
  AOI22_X1 U165 ( .A1(H[63]), .A2(n1441), .B1(G[63]), .B2(n1435), .ZN(n30) );
  AOI22_X1 U166 ( .A1(F[39]), .A2(n1427), .B1(E[39]), .B2(n1421), .ZN(n137) );
  NAND4_X1 U167 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(Y[39]) );
  AOI22_X1 U168 ( .A1(B[39]), .A2(n1403), .B1(A[39]), .B2(n1397), .ZN(n135) );
  AOI22_X1 U169 ( .A1(D[39]), .A2(n1415), .B1(C[39]), .B2(n1409), .ZN(n136) );
  AOI22_X1 U170 ( .A1(H[39]), .A2(n1439), .B1(G[39]), .B2(n1433), .ZN(n138) );
  AOI22_X1 U171 ( .A1(F[30]), .A2(n1426), .B1(E[30]), .B2(n1420), .ZN(n173) );
  AOI22_X1 U172 ( .A1(F[37]), .A2(n1427), .B1(E[37]), .B2(n1421), .ZN(n145) );
  AOI22_X1 U173 ( .A1(F[35]), .A2(n1427), .B1(E[35]), .B2(n1421), .ZN(n153) );
  AOI22_X1 U174 ( .A1(F[38]), .A2(n1427), .B1(E[38]), .B2(n1421), .ZN(n141) );
  AOI22_X1 U175 ( .A1(D[31]), .A2(n1415), .B1(C[31]), .B2(n1409), .ZN(n168) );
  AOI22_X1 U176 ( .A1(D[33]), .A2(n1415), .B1(C[33]), .B2(n1409), .ZN(n160) );
  AOI22_X1 U177 ( .A1(D[34]), .A2(n1415), .B1(C[34]), .B2(n1409), .ZN(n156) );
  AOI22_X1 U178 ( .A1(D[32]), .A2(n1415), .B1(C[32]), .B2(n1409), .ZN(n164) );
  NAND4_X1 U179 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(Y[35]) );
  AOI22_X1 U180 ( .A1(B[35]), .A2(n1403), .B1(A[35]), .B2(n1397), .ZN(n151) );
  AOI22_X1 U181 ( .A1(H[35]), .A2(n1439), .B1(G[35]), .B2(n1433), .ZN(n154) );
  AOI22_X1 U182 ( .A1(D[35]), .A2(n1415), .B1(C[35]), .B2(n1409), .ZN(n152) );
  NAND4_X1 U183 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(Y[30]) );
  AOI22_X1 U184 ( .A1(D[30]), .A2(n1414), .B1(C[30]), .B2(n1408), .ZN(n172) );
  AOI22_X1 U185 ( .A1(H[30]), .A2(n1438), .B1(G[30]), .B2(n1432), .ZN(n174) );
  AOI22_X1 U186 ( .A1(B[30]), .A2(n1402), .B1(A[30]), .B2(n1396), .ZN(n171) );
  NAND4_X1 U187 ( .A1(n143), .A2(n144), .A3(n145), .A4(n146), .ZN(Y[37]) );
  AOI22_X1 U188 ( .A1(B[37]), .A2(n1403), .B1(A[37]), .B2(n1397), .ZN(n143) );
  AOI22_X1 U189 ( .A1(H[37]), .A2(n1439), .B1(G[37]), .B2(n1433), .ZN(n146) );
  AOI22_X1 U190 ( .A1(D[37]), .A2(n1415), .B1(C[37]), .B2(n1409), .ZN(n144) );
  NAND4_X1 U191 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .ZN(Y[38]) );
  AOI22_X1 U192 ( .A1(B[38]), .A2(n1403), .B1(A[38]), .B2(n1397), .ZN(n139) );
  AOI22_X1 U193 ( .A1(H[38]), .A2(n1439), .B1(G[38]), .B2(n1433), .ZN(n142) );
  AOI22_X1 U194 ( .A1(D[38]), .A2(n1415), .B1(C[38]), .B2(n1409), .ZN(n140) );
  NAND4_X1 U195 ( .A1(n127), .A2(n128), .A3(n129), .A4(n130), .ZN(Y[40]) );
  AOI22_X1 U196 ( .A1(B[40]), .A2(n1403), .B1(A[40]), .B2(n1397), .ZN(n127) );
  AOI22_X1 U197 ( .A1(D[40]), .A2(n1415), .B1(C[40]), .B2(n1409), .ZN(n128) );
  AOI22_X1 U198 ( .A1(H[40]), .A2(n1439), .B1(G[40]), .B2(n1433), .ZN(n130) );
  NAND4_X1 U199 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U200 ( .A1(H[31]), .A2(n1439), .B1(G[31]), .B2(n1433), .ZN(n170) );
  AOI22_X1 U201 ( .A1(B[31]), .A2(n1403), .B1(A[31]), .B2(n1397), .ZN(n167) );
  AOI22_X1 U202 ( .A1(F[31]), .A2(n1427), .B1(E[31]), .B2(n1421), .ZN(n169) );
  NAND4_X1 U203 ( .A1(n147), .A2(n148), .A3(n149), .A4(n150), .ZN(Y[36]) );
  AOI22_X1 U204 ( .A1(H[36]), .A2(n1439), .B1(G[36]), .B2(n1433), .ZN(n150) );
  AOI22_X1 U205 ( .A1(B[36]), .A2(n1403), .B1(A[36]), .B2(n1397), .ZN(n147) );
  AOI22_X1 U206 ( .A1(D[36]), .A2(n1415), .B1(C[36]), .B2(n1409), .ZN(n148) );
  NAND4_X1 U207 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(Y[33]) );
  AOI22_X1 U208 ( .A1(B[33]), .A2(n1403), .B1(A[33]), .B2(n1397), .ZN(n159) );
  AOI22_X1 U209 ( .A1(H[33]), .A2(n1439), .B1(G[33]), .B2(n1433), .ZN(n162) );
  AOI22_X1 U210 ( .A1(F[33]), .A2(n1427), .B1(E[33]), .B2(n1421), .ZN(n161) );
  NAND4_X1 U211 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .ZN(Y[34]) );
  AOI22_X1 U212 ( .A1(B[34]), .A2(n1403), .B1(A[34]), .B2(n1397), .ZN(n155) );
  AOI22_X1 U213 ( .A1(H[34]), .A2(n1439), .B1(G[34]), .B2(n1433), .ZN(n158) );
  AOI22_X1 U214 ( .A1(F[34]), .A2(n1427), .B1(E[34]), .B2(n1421), .ZN(n157) );
  NAND4_X1 U215 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .ZN(Y[32]) );
  AOI22_X1 U216 ( .A1(B[32]), .A2(n1403), .B1(A[32]), .B2(n1397), .ZN(n163) );
  AOI22_X1 U217 ( .A1(H[32]), .A2(n1439), .B1(G[32]), .B2(n1433), .ZN(n166) );
  AOI22_X1 U218 ( .A1(F[32]), .A2(n1427), .B1(E[32]), .B2(n1421), .ZN(n165) );
  AOI22_X1 U219 ( .A1(F[40]), .A2(n1427), .B1(E[40]), .B2(n1421), .ZN(n129) );
  AOI22_X1 U220 ( .A1(F[36]), .A2(n1427), .B1(E[36]), .B2(n1421), .ZN(n149) );
  NAND4_X1 U221 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(Y[0]) );
  AOI22_X1 U222 ( .A1(B[0]), .A2(n1401), .B1(A[0]), .B2(n1395), .ZN(n263) );
  AOI22_X1 U223 ( .A1(D[0]), .A2(n1413), .B1(C[0]), .B2(n1407), .ZN(n264) );
  AOI22_X1 U224 ( .A1(F[0]), .A2(n1425), .B1(E[0]), .B2(n1419), .ZN(n265) );
  AOI22_X1 U225 ( .A1(H[7]), .A2(n1442), .B1(G[7]), .B2(n1436), .ZN(n22) );
  AOI22_X1 U226 ( .A1(H[11]), .A2(n1437), .B1(G[11]), .B2(n1431), .ZN(n258) );
  AOI22_X1 U227 ( .A1(H[15]), .A2(n1437), .B1(G[15]), .B2(n1431), .ZN(n242) );
  AOI22_X1 U228 ( .A1(H[23]), .A2(n1438), .B1(G[23]), .B2(n1432), .ZN(n206) );
  AOI22_X1 U229 ( .A1(H[27]), .A2(n1438), .B1(G[27]), .B2(n1432), .ZN(n190) );
  AOI22_X1 U230 ( .A1(H[19]), .A2(n1437), .B1(G[19]), .B2(n1431), .ZN(n226) );
  AOI22_X1 U231 ( .A1(H[21]), .A2(n1438), .B1(G[21]), .B2(n1432), .ZN(n214) );
  AOI22_X1 U232 ( .A1(H[29]), .A2(n1438), .B1(G[29]), .B2(n1432), .ZN(n182) );
  AOI22_X1 U233 ( .A1(H[5]), .A2(n1441), .B1(G[5]), .B2(n1435), .ZN(n46) );
  AOI22_X1 U234 ( .A1(H[9]), .A2(n1442), .B1(G[9]), .B2(n1436), .ZN(n6) );
  AOI22_X1 U235 ( .A1(H[13]), .A2(n1437), .B1(G[13]), .B2(n1431), .ZN(n250) );
  AOI22_X1 U236 ( .A1(H[17]), .A2(n1437), .B1(G[17]), .B2(n1431), .ZN(n234) );
  AOI22_X1 U237 ( .A1(H[25]), .A2(n1438), .B1(G[25]), .B2(n1432), .ZN(n198) );
  AOI22_X1 U238 ( .A1(H[3]), .A2(n1439), .B1(G[3]), .B2(n1433), .ZN(n134) );
  AOI22_X1 U239 ( .A1(H[4]), .A2(n1440), .B1(G[4]), .B2(n1434), .ZN(n90) );
  AOI22_X1 U240 ( .A1(H[8]), .A2(n1442), .B1(G[8]), .B2(n1436), .ZN(n18) );
  AOI22_X1 U241 ( .A1(H[12]), .A2(n1437), .B1(G[12]), .B2(n1431), .ZN(n254) );
  AOI22_X1 U242 ( .A1(H[16]), .A2(n1437), .B1(G[16]), .B2(n1431), .ZN(n238) );
  AOI22_X1 U243 ( .A1(H[20]), .A2(n1438), .B1(G[20]), .B2(n1432), .ZN(n218) );
  AOI22_X1 U244 ( .A1(H[24]), .A2(n1438), .B1(G[24]), .B2(n1432), .ZN(n202) );
  AOI22_X1 U245 ( .A1(H[28]), .A2(n1438), .B1(G[28]), .B2(n1432), .ZN(n186) );
  AOI22_X1 U246 ( .A1(H[6]), .A2(n1442), .B1(G[6]), .B2(n1436), .ZN(n26) );
  AOI22_X1 U247 ( .A1(H[10]), .A2(n1437), .B1(G[10]), .B2(n1431), .ZN(n262) );
  AOI22_X1 U248 ( .A1(H[14]), .A2(n1437), .B1(G[14]), .B2(n1431), .ZN(n246) );
  AOI22_X1 U249 ( .A1(H[18]), .A2(n1437), .B1(G[18]), .B2(n1431), .ZN(n230) );
  AOI22_X1 U250 ( .A1(H[22]), .A2(n1438), .B1(G[22]), .B2(n1432), .ZN(n210) );
  AOI22_X1 U251 ( .A1(H[26]), .A2(n1438), .B1(G[26]), .B2(n1432), .ZN(n194) );
  AOI22_X1 U252 ( .A1(H[2]), .A2(n1438), .B1(G[2]), .B2(n1432), .ZN(n178) );
  AOI22_X1 U253 ( .A1(H[1]), .A2(n1437), .B1(G[1]), .B2(n1431), .ZN(n222) );
  NAND4_X1 U254 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(Y[15]) );
  AOI22_X1 U255 ( .A1(B[15]), .A2(n1401), .B1(A[15]), .B2(n1395), .ZN(n239) );
  AOI22_X1 U256 ( .A1(D[15]), .A2(n1413), .B1(C[15]), .B2(n1407), .ZN(n240) );
  AOI22_X1 U257 ( .A1(F[15]), .A2(n1425), .B1(E[15]), .B2(n1419), .ZN(n241) );
  NAND4_X1 U258 ( .A1(n203), .A2(n204), .A3(n205), .A4(n206), .ZN(Y[23]) );
  AOI22_X1 U259 ( .A1(B[23]), .A2(n1402), .B1(A[23]), .B2(n1396), .ZN(n203) );
  AOI22_X1 U260 ( .A1(D[23]), .A2(n1414), .B1(C[23]), .B2(n1408), .ZN(n204) );
  AOI22_X1 U261 ( .A1(F[23]), .A2(n1426), .B1(E[23]), .B2(n1420), .ZN(n205) );
  NAND4_X1 U262 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(Y[27]) );
  AOI22_X1 U263 ( .A1(B[27]), .A2(n1402), .B1(A[27]), .B2(n1396), .ZN(n187) );
  AOI22_X1 U264 ( .A1(D[27]), .A2(n1414), .B1(C[27]), .B2(n1408), .ZN(n188) );
  AOI22_X1 U265 ( .A1(F[27]), .A2(n1426), .B1(E[27]), .B2(n1420), .ZN(n189) );
  NAND4_X1 U266 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(Y[19]) );
  AOI22_X1 U267 ( .A1(B[19]), .A2(n1401), .B1(A[19]), .B2(n1395), .ZN(n223) );
  AOI22_X1 U268 ( .A1(D[19]), .A2(n1413), .B1(C[19]), .B2(n1407), .ZN(n224) );
  AOI22_X1 U269 ( .A1(F[19]), .A2(n1425), .B1(E[19]), .B2(n1419), .ZN(n225) );
  NAND4_X1 U270 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(Y[21]) );
  AOI22_X1 U271 ( .A1(B[21]), .A2(n1402), .B1(A[21]), .B2(n1396), .ZN(n211) );
  AOI22_X1 U272 ( .A1(D[21]), .A2(n1414), .B1(C[21]), .B2(n1408), .ZN(n212) );
  AOI22_X1 U273 ( .A1(F[21]), .A2(n1426), .B1(E[21]), .B2(n1420), .ZN(n213) );
  NAND4_X1 U274 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(Y[29]) );
  AOI22_X1 U275 ( .A1(B[29]), .A2(n1402), .B1(A[29]), .B2(n1396), .ZN(n179) );
  AOI22_X1 U276 ( .A1(D[29]), .A2(n1414), .B1(C[29]), .B2(n1408), .ZN(n180) );
  AOI22_X1 U277 ( .A1(F[29]), .A2(n1426), .B1(E[29]), .B2(n1420), .ZN(n181) );
  NAND4_X1 U278 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(Y[5]) );
  AOI22_X1 U279 ( .A1(B[5]), .A2(n1405), .B1(A[5]), .B2(n1399), .ZN(n43) );
  AOI22_X1 U280 ( .A1(D[5]), .A2(n1417), .B1(C[5]), .B2(n1411), .ZN(n44) );
  AOI22_X1 U281 ( .A1(F[5]), .A2(n1429), .B1(E[5]), .B2(n1423), .ZN(n45) );
  NAND4_X1 U282 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(Y[9]) );
  AOI22_X1 U283 ( .A1(B[9]), .A2(n1406), .B1(A[9]), .B2(n1400), .ZN(n3) );
  AOI22_X1 U284 ( .A1(D[9]), .A2(n1418), .B1(C[9]), .B2(n1412), .ZN(n4) );
  AOI22_X1 U285 ( .A1(F[9]), .A2(n1430), .B1(E[9]), .B2(n1424), .ZN(n5) );
  NAND4_X1 U286 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(Y[17]) );
  AOI22_X1 U287 ( .A1(B[17]), .A2(n1401), .B1(A[17]), .B2(n1395), .ZN(n231) );
  AOI22_X1 U288 ( .A1(D[17]), .A2(n1413), .B1(C[17]), .B2(n1407), .ZN(n232) );
  AOI22_X1 U289 ( .A1(F[17]), .A2(n1425), .B1(E[17]), .B2(n1419), .ZN(n233) );
  NAND4_X1 U290 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(Y[3]) );
  AOI22_X1 U291 ( .A1(B[3]), .A2(n1403), .B1(A[3]), .B2(n1397), .ZN(n131) );
  AOI22_X1 U292 ( .A1(D[3]), .A2(n1415), .B1(C[3]), .B2(n1409), .ZN(n132) );
  AOI22_X1 U293 ( .A1(F[3]), .A2(n1427), .B1(E[3]), .B2(n1421), .ZN(n133) );
  NAND4_X1 U294 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(Y[7]) );
  AOI22_X1 U295 ( .A1(B[7]), .A2(n1406), .B1(A[7]), .B2(n1400), .ZN(n19) );
  AOI22_X1 U296 ( .A1(D[7]), .A2(n1418), .B1(C[7]), .B2(n1412), .ZN(n20) );
  AOI22_X1 U297 ( .A1(F[7]), .A2(n1430), .B1(E[7]), .B2(n1424), .ZN(n21) );
  NAND4_X1 U298 ( .A1(n255), .A2(n256), .A3(n257), .A4(n258), .ZN(Y[11]) );
  AOI22_X1 U299 ( .A1(B[11]), .A2(n1401), .B1(A[11]), .B2(n1395), .ZN(n255) );
  AOI22_X1 U300 ( .A1(D[11]), .A2(n1413), .B1(C[11]), .B2(n1407), .ZN(n256) );
  AOI22_X1 U301 ( .A1(F[11]), .A2(n1425), .B1(E[11]), .B2(n1419), .ZN(n257) );
  NAND4_X1 U302 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(Y[13]) );
  AOI22_X1 U303 ( .A1(B[13]), .A2(n1401), .B1(A[13]), .B2(n1395), .ZN(n247) );
  AOI22_X1 U304 ( .A1(D[13]), .A2(n1413), .B1(C[13]), .B2(n1407), .ZN(n248) );
  AOI22_X1 U305 ( .A1(F[13]), .A2(n1425), .B1(E[13]), .B2(n1419), .ZN(n249) );
  NAND4_X1 U306 ( .A1(n195), .A2(n196), .A3(n197), .A4(n198), .ZN(Y[25]) );
  AOI22_X1 U307 ( .A1(B[25]), .A2(n1402), .B1(A[25]), .B2(n1396), .ZN(n195) );
  AOI22_X1 U308 ( .A1(D[25]), .A2(n1414), .B1(C[25]), .B2(n1408), .ZN(n196) );
  AOI22_X1 U309 ( .A1(F[25]), .A2(n1426), .B1(E[25]), .B2(n1420), .ZN(n197) );
  NAND4_X1 U310 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .ZN(Y[4]) );
  AOI22_X1 U311 ( .A1(B[4]), .A2(n1404), .B1(A[4]), .B2(n1398), .ZN(n87) );
  AOI22_X1 U312 ( .A1(D[4]), .A2(n1416), .B1(C[4]), .B2(n1410), .ZN(n88) );
  AOI22_X1 U313 ( .A1(F[4]), .A2(n1428), .B1(E[4]), .B2(n1422), .ZN(n89) );
  NAND4_X1 U314 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(Y[6]) );
  AOI22_X1 U315 ( .A1(B[6]), .A2(n1406), .B1(A[6]), .B2(n1400), .ZN(n23) );
  AOI22_X1 U316 ( .A1(D[6]), .A2(n1418), .B1(C[6]), .B2(n1412), .ZN(n24) );
  AOI22_X1 U317 ( .A1(F[6]), .A2(n1430), .B1(E[6]), .B2(n1424), .ZN(n25) );
  NAND4_X1 U318 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(Y[8]) );
  AOI22_X1 U319 ( .A1(B[8]), .A2(n1406), .B1(A[8]), .B2(n1400), .ZN(n15) );
  AOI22_X1 U320 ( .A1(D[8]), .A2(n1418), .B1(C[8]), .B2(n1412), .ZN(n16) );
  AOI22_X1 U321 ( .A1(F[8]), .A2(n1430), .B1(E[8]), .B2(n1424), .ZN(n17) );
  NAND4_X1 U322 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(Y[10]) );
  AOI22_X1 U323 ( .A1(B[10]), .A2(n1401), .B1(A[10]), .B2(n1395), .ZN(n259) );
  AOI22_X1 U324 ( .A1(D[10]), .A2(n1413), .B1(C[10]), .B2(n1407), .ZN(n260) );
  AOI22_X1 U325 ( .A1(F[10]), .A2(n1425), .B1(E[10]), .B2(n1419), .ZN(n261) );
  NAND4_X1 U326 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(Y[12]) );
  AOI22_X1 U327 ( .A1(B[12]), .A2(n1401), .B1(A[12]), .B2(n1395), .ZN(n251) );
  AOI22_X1 U328 ( .A1(D[12]), .A2(n1413), .B1(C[12]), .B2(n1407), .ZN(n252) );
  AOI22_X1 U329 ( .A1(F[12]), .A2(n1425), .B1(E[12]), .B2(n1419), .ZN(n253) );
  NAND4_X1 U330 ( .A1(n243), .A2(n244), .A3(n245), .A4(n246), .ZN(Y[14]) );
  AOI22_X1 U331 ( .A1(B[14]), .A2(n1401), .B1(A[14]), .B2(n1395), .ZN(n243) );
  AOI22_X1 U332 ( .A1(D[14]), .A2(n1413), .B1(C[14]), .B2(n1407), .ZN(n244) );
  AOI22_X1 U333 ( .A1(F[14]), .A2(n1425), .B1(E[14]), .B2(n1419), .ZN(n245) );
  NAND4_X1 U334 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(Y[16]) );
  AOI22_X1 U335 ( .A1(B[16]), .A2(n1401), .B1(A[16]), .B2(n1395), .ZN(n235) );
  AOI22_X1 U336 ( .A1(D[16]), .A2(n1413), .B1(C[16]), .B2(n1407), .ZN(n236) );
  AOI22_X1 U337 ( .A1(F[16]), .A2(n1425), .B1(E[16]), .B2(n1419), .ZN(n237) );
  NAND4_X1 U338 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(Y[18]) );
  AOI22_X1 U339 ( .A1(B[18]), .A2(n1401), .B1(A[18]), .B2(n1395), .ZN(n227) );
  AOI22_X1 U340 ( .A1(D[18]), .A2(n1413), .B1(C[18]), .B2(n1407), .ZN(n228) );
  AOI22_X1 U341 ( .A1(F[18]), .A2(n1425), .B1(E[18]), .B2(n1419), .ZN(n229) );
  NAND4_X1 U342 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(Y[20]) );
  AOI22_X1 U343 ( .A1(B[20]), .A2(n1402), .B1(A[20]), .B2(n1396), .ZN(n215) );
  AOI22_X1 U344 ( .A1(D[20]), .A2(n1414), .B1(C[20]), .B2(n1408), .ZN(n216) );
  AOI22_X1 U345 ( .A1(F[20]), .A2(n1426), .B1(E[20]), .B2(n1420), .ZN(n217) );
  NAND4_X1 U346 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(Y[22]) );
  AOI22_X1 U347 ( .A1(B[22]), .A2(n1402), .B1(A[22]), .B2(n1396), .ZN(n207) );
  AOI22_X1 U348 ( .A1(D[22]), .A2(n1414), .B1(C[22]), .B2(n1408), .ZN(n208) );
  AOI22_X1 U349 ( .A1(F[22]), .A2(n1426), .B1(E[22]), .B2(n1420), .ZN(n209) );
  NAND4_X1 U350 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(Y[24]) );
  AOI22_X1 U351 ( .A1(B[24]), .A2(n1402), .B1(A[24]), .B2(n1396), .ZN(n199) );
  AOI22_X1 U352 ( .A1(D[24]), .A2(n1414), .B1(C[24]), .B2(n1408), .ZN(n200) );
  AOI22_X1 U353 ( .A1(F[24]), .A2(n1426), .B1(E[24]), .B2(n1420), .ZN(n201) );
  NAND4_X1 U354 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(Y[26]) );
  AOI22_X1 U355 ( .A1(B[26]), .A2(n1402), .B1(A[26]), .B2(n1396), .ZN(n191) );
  AOI22_X1 U356 ( .A1(D[26]), .A2(n1414), .B1(C[26]), .B2(n1408), .ZN(n192) );
  AOI22_X1 U357 ( .A1(F[26]), .A2(n1426), .B1(E[26]), .B2(n1420), .ZN(n193) );
  NAND4_X1 U358 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(Y[28]) );
  AOI22_X1 U359 ( .A1(B[28]), .A2(n1402), .B1(A[28]), .B2(n1396), .ZN(n183) );
  AOI22_X1 U360 ( .A1(D[28]), .A2(n1414), .B1(C[28]), .B2(n1408), .ZN(n184) );
  AOI22_X1 U361 ( .A1(F[28]), .A2(n1426), .B1(E[28]), .B2(n1420), .ZN(n185) );
  NAND4_X1 U362 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(Y[2]) );
  AOI22_X1 U363 ( .A1(B[2]), .A2(n1402), .B1(A[2]), .B2(n1396), .ZN(n175) );
  AOI22_X1 U364 ( .A1(D[2]), .A2(n1414), .B1(C[2]), .B2(n1408), .ZN(n176) );
  AOI22_X1 U365 ( .A1(F[2]), .A2(n1426), .B1(E[2]), .B2(n1420), .ZN(n177) );
  NAND4_X1 U366 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(Y[1]) );
  AOI22_X1 U367 ( .A1(B[1]), .A2(n1401), .B1(A[1]), .B2(n1395), .ZN(n219) );
  AOI22_X1 U368 ( .A1(D[1]), .A2(n1413), .B1(C[1]), .B2(n1407), .ZN(n220) );
  AOI22_X1 U369 ( .A1(F[1]), .A2(n1425), .B1(E[1]), .B2(n1419), .ZN(n221) );
  AOI22_X1 U370 ( .A1(H[0]), .A2(n1437), .B1(G[0]), .B2(n1431), .ZN(n266) );
  CLKBUF_X1 U371 ( .A(n14), .Z(n1400) );
  CLKBUF_X1 U372 ( .A(n13), .Z(n1406) );
  CLKBUF_X1 U373 ( .A(n12), .Z(n1412) );
  CLKBUF_X1 U374 ( .A(n11), .Z(n1418) );
  CLKBUF_X1 U375 ( .A(n10), .Z(n1424) );
  CLKBUF_X1 U376 ( .A(n9), .Z(n1430) );
  CLKBUF_X1 U377 ( .A(n8), .Z(n1436) );
  CLKBUF_X1 U378 ( .A(n7), .Z(n1442) );
endmodule


module RCA_NBIT64_0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net513018, net513010, net513005, net513004, net513003, net513001,
         net512989, net512987, net512986, net512977, net512976, net512975,
         net512964, net512962, net512961, net512958, net512956, net512953,
         net512943, net512908, net512907, net512906, net512905, net512903,
         net512901, net512900, net512899, net512889, net512883, net512825,
         net512809, net512807, net512806, net512804, net537302, net537536,
         net537535, net537976, net538262, net538396, net512944, net512942,
         net512938, net512876, net512875, net512868, net512864, net512863,
         net512862, net512861, net512990, net512827, net512808, net512881,
         net512869, net512867, net512866, net537046, net512870, net512871,
         net512829, net512810, net512937, net512936, net512935, net512934, n2,
         n3, n4, n6, n7, n8, n9, n10, n11, n12, n16, n17, n18, n19, n21, n23,
         n25, n29, n30, n31, n32, n33, n34, n35, n38, n39, n41, n42, n43, n44,
         n45, n47, n51, n52, n53, n54, n56, n58, n59, n60, n62, n64, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n77, n80, n81, n82, n84, n85, n87,
         n89, n90, n91, n92, n94, n95, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n123, n124, n126, n127, n128,
         n129, n130, n131, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n151, n152, n153,
         n155, n156, n157, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n174, n176, n177, n179, n180, n181,
         n183, n184, n185, n187, n188, n189, n192, n193, n194, n195, n196,
         n197, n198, n200, n202, n203, n205, n206, n207, n209, n210, n211,
         n213, n214, n215, n218, n219, n220, n221, n222, n223, n224, n226,
         n228, n229, n230, n231, n233, n234, n235, n237, n238, n239, n240,
         n242, n243, n244, n246, n247, n248, n249, n251, n252, n253, n254,
         n256, n257, n259, n260, n261, n262, n263, n264, n265, n266, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n292,
         n293, n294, n295, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n312, n313, n314, n315, n316, n317,
         n318, n321, n322, n324, n325, n326, n327, n328, n329, n331, n332,
         n333, n335, n336, n337, n338, n339, n340, n341, n342, n344, n345,
         n347, n348, n349, n350, n351, n353, n354, n355, n356, n357, n359,
         n360, n361, n362, n363, n364, n365, n366, n369, n372, n373, n374,
         n375, n377, n379, n380, n381, n382, n383, n384, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n400, n401,
         n402, n403, n405, n406, n407, n408, n411, n412, n413, n414, n415,
         n416, n417, n423, n424, n425, n426, n427, n428, n429, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555;

  NAND3_X1 U78 ( .A1(net512975), .A2(net512976), .A3(net512977), .ZN(n34) );
  NAND3_X1 U91 ( .A1(net538396), .A2(n492), .A3(net512989), .ZN(net513010) );
  OR2_X2 U159 ( .A1(A[5]), .A2(B[5]), .ZN(n116) );
  NAND3_X1 U506 ( .A1(n91), .A2(n8), .A3(n92), .ZN(n89) );
  NAND3_X1 U562 ( .A1(net512806), .A2(n488), .A3(net512804), .ZN(n349) );
  NAND3_X1 U575 ( .A1(n59), .A2(n439), .A3(n393), .ZN(net512976) );
  NAND3_X1 U576 ( .A1(n454), .A2(n106), .A3(n108), .ZN(n393) );
  NAND3_X1 U577 ( .A1(net513010), .A2(n397), .A3(net513005), .ZN(n395) );
  NAND3_X1 U583 ( .A1(n439), .A2(n67), .A3(n230), .ZN(n417) );
  NAND3_X1 U587 ( .A1(n91), .A2(n8), .A3(n92), .ZN(n108) );
  NAND3_X1 U589 ( .A1(n116), .A2(A[4]), .A3(n436), .ZN(n424) );
  OR2_X1 U2 ( .A1(B[11]), .A2(A[11]), .ZN(n407) );
  AND2_X1 U3 ( .A1(n429), .A2(n390), .ZN(SUM[0]) );
  OR2_X1 U4 ( .A1(B[16]), .A2(A[16]), .ZN(net512943) );
  OR2_X1 U5 ( .A1(B[26]), .A2(A[26]), .ZN(net512868) );
  AND2_X1 U6 ( .A1(n364), .A2(n363), .ZN(n432) );
  OAI21_X2 U7 ( .B1(n9), .B2(n31), .A(net512899), .ZN(net512829) );
  CLKBUF_X1 U8 ( .A(A[11]), .Z(n433) );
  CLKBUF_X1 U9 ( .A(net512827), .Z(n434) );
  OAI21_X1 U10 ( .B1(n474), .B2(net512810), .A(net512829), .ZN(n435) );
  BUF_X1 U11 ( .A(B[4]), .Z(n436) );
  BUF_X1 U12 ( .A(A[2]), .Z(n437) );
  OR2_X1 U13 ( .A1(B[3]), .A2(A[3]), .ZN(n438) );
  OR2_X1 U14 ( .A1(B[3]), .A2(A[3]), .ZN(n169) );
  AND4_X1 U15 ( .A1(n109), .A2(n116), .A3(n123), .A4(n102), .ZN(n439) );
  OR2_X2 U16 ( .A1(B[14]), .A2(A[14]), .ZN(net512989) );
  AND2_X1 U17 ( .A1(n82), .A2(n60), .ZN(n440) );
  AND2_X2 U18 ( .A1(n53), .A2(n440), .ZN(n59) );
  OR2_X2 U19 ( .A1(B[9]), .A2(A[9]), .ZN(n411) );
  CLKBUF_X1 U20 ( .A(n394), .Z(n442) );
  XOR2_X1 U21 ( .A(n19), .B(n441), .Z(SUM[12]) );
  NAND2_X1 U22 ( .A1(n403), .A2(net512977), .ZN(n441) );
  NAND4_X1 U23 ( .A1(n109), .A2(n116), .A3(n123), .A4(n102), .ZN(n394) );
  OR2_X1 U24 ( .A1(B[17]), .A2(A[17]), .ZN(net512944) );
  AND2_X1 U25 ( .A1(n415), .A2(n80), .ZN(n443) );
  AND3_X1 U26 ( .A1(n417), .A2(n416), .A3(n443), .ZN(n68) );
  INV_X1 U27 ( .A(n230), .ZN(n444) );
  AND2_X1 U28 ( .A1(n379), .A2(n359), .ZN(n445) );
  AND2_X1 U29 ( .A1(n379), .A2(n359), .ZN(n54) );
  XNOR2_X1 U30 ( .A(n446), .B(n447), .ZN(SUM[19]) );
  NAND2_X1 U31 ( .A1(n23), .A2(net512942), .ZN(n446) );
  NAND2_X1 U32 ( .A1(net512935), .A2(net512937), .ZN(n447) );
  AND3_X1 U33 ( .A1(net512977), .A2(net512976), .A3(net512975), .ZN(n448) );
  AND3_X1 U34 ( .A1(net512975), .A2(net512976), .A3(net512977), .ZN(net538262)
         );
  OR2_X1 U35 ( .A1(A[4]), .A2(B[4]), .ZN(n449) );
  OR2_X1 U36 ( .A1(A[4]), .A2(n436), .ZN(n123) );
  INV_X1 U37 ( .A(n45), .ZN(n450) );
  AOI21_X1 U38 ( .B1(n435), .B2(net512871), .A(n542), .ZN(n451) );
  XNOR2_X1 U39 ( .A(n29), .B(n452), .ZN(SUM[14]) );
  AND2_X1 U40 ( .A1(net512989), .A2(net513005), .ZN(n452) );
  NAND3_X1 U41 ( .A1(n169), .A2(B[2]), .A3(A[2]), .ZN(n453) );
  NAND3_X1 U42 ( .A1(n438), .A2(B[2]), .A3(n437), .ZN(n454) );
  NAND3_X1 U43 ( .A1(n169), .A2(B[2]), .A3(A[2]), .ZN(n90) );
  OR2_X2 U44 ( .A1(n256), .A2(n69), .ZN(n324) );
  NAND3_X1 U45 ( .A1(n356), .A2(n355), .A3(n432), .ZN(net512807) );
  OR2_X1 U46 ( .A1(B[30]), .A2(A[30]), .ZN(n355) );
  NAND2_X1 U47 ( .A1(n348), .A2(n458), .ZN(n455) );
  AND2_X1 U48 ( .A1(n455), .A2(n456), .ZN(n344) );
  OR2_X1 U49 ( .A1(n457), .A2(n326), .ZN(n456) );
  INV_X1 U50 ( .A(n335), .ZN(n457) );
  AND2_X1 U51 ( .A1(n349), .A2(n335), .ZN(n458) );
  AND2_X1 U52 ( .A1(n41), .A2(net512989), .ZN(n38) );
  OR2_X2 U53 ( .A1(B[6]), .A2(A[6]), .ZN(n102) );
  XNOR2_X1 U54 ( .A(n488), .B(n459), .ZN(SUM[16]) );
  NAND2_X1 U55 ( .A1(net512943), .A2(n42), .ZN(n459) );
  XOR2_X1 U56 ( .A(n435), .B(n460), .Z(SUM[24]) );
  AND2_X1 U57 ( .A1(net512871), .A2(net512870), .ZN(n460) );
  XOR2_X1 U58 ( .A(n461), .B(n97), .Z(SUM[7]) );
  AND2_X1 U59 ( .A1(n109), .A2(n110), .ZN(n461) );
  XOR2_X1 U60 ( .A(n52), .B(n462), .Z(SUM[30]) );
  AND2_X1 U61 ( .A1(n355), .A2(n361), .ZN(n462) );
  XNOR2_X1 U62 ( .A(n463), .B(n56), .ZN(SUM[10]) );
  AND4_X1 U63 ( .A1(n80), .A2(n415), .A3(n416), .A4(n417), .ZN(n463) );
  XOR2_X1 U64 ( .A(n467), .B(n464), .Z(SUM[21]) );
  NAND2_X1 U65 ( .A1(n387), .A2(net512907), .ZN(n464) );
  INV_X1 U66 ( .A(n233), .ZN(n481) );
  INV_X1 U67 ( .A(n7), .ZN(n488) );
  OAI211_X1 U68 ( .C1(n235), .C2(n482), .A(n237), .B(n238), .ZN(n233) );
  AOI21_X1 U69 ( .B1(n239), .B2(n240), .A(n524), .ZN(n238) );
  INV_X1 U70 ( .A(n435), .ZN(n472) );
  OAI21_X1 U71 ( .B1(n7), .B2(net512808), .A(n495), .ZN(net537976) );
  AOI21_X1 U72 ( .B1(n501), .B2(n434), .A(n499), .ZN(n362) );
  INV_X1 U73 ( .A(net512810), .ZN(n501) );
  INV_X1 U74 ( .A(n33), .ZN(n474) );
  OAI21_X1 U75 ( .B1(n6), .B2(net512808), .A(n495), .ZN(n33) );
  AND2_X1 U76 ( .A1(n21), .A2(n35), .ZN(n6) );
  OAI21_X1 U77 ( .B1(n249), .B2(n520), .A(n72), .ZN(n237) );
  INV_X1 U79 ( .A(n251), .ZN(n520) );
  NAND2_X1 U80 ( .A1(n273), .A2(n251), .ZN(n271) );
  NAND2_X1 U81 ( .A1(n108), .A2(n62), .ZN(n230) );
  INV_X1 U82 ( .A(net512827), .ZN(n495) );
  AND2_X1 U83 ( .A1(n21), .A2(n35), .ZN(n7) );
  INV_X1 U84 ( .A(n205), .ZN(n480) );
  INV_X1 U85 ( .A(n179), .ZN(n479) );
  INV_X1 U86 ( .A(n261), .ZN(n518) );
  INV_X1 U87 ( .A(n103), .ZN(n491) );
  INV_X1 U88 ( .A(n147), .ZN(n477) );
  NAND2_X1 U89 ( .A1(n2), .A2(n59), .ZN(net512975) );
  OR2_X1 U90 ( .A1(n94), .A2(n490), .ZN(n2) );
  NAND2_X1 U92 ( .A1(n34), .A2(n25), .ZN(n35) );
  NAND2_X1 U93 ( .A1(n104), .A2(n103), .ZN(n101) );
  NAND2_X1 U94 ( .A1(n64), .A2(n51), .ZN(n416) );
  NOR2_X1 U95 ( .A1(n119), .A2(n120), .ZN(n113) );
  NAND2_X1 U96 ( .A1(n491), .A2(n8), .ZN(n120) );
  NAND2_X1 U97 ( .A1(n91), .A2(n92), .ZN(n119) );
  NOR2_X1 U98 ( .A1(n124), .A2(n537), .ZN(SUM[64]) );
  INV_X1 U99 ( .A(n313), .ZN(n551) );
  XNOR2_X1 U100 ( .A(n58), .B(n465), .ZN(SUM[8]) );
  NAND2_X1 U101 ( .A1(n428), .A2(n82), .ZN(n465) );
  NOR2_X1 U102 ( .A1(n544), .A2(n545), .ZN(n77) );
  INV_X1 U103 ( .A(n80), .ZN(n544) );
  NAND2_X1 U104 ( .A1(n492), .A2(net513004), .ZN(net513018) );
  OAI211_X1 U105 ( .C1(n498), .C2(n42), .A(n43), .B(net512942), .ZN(net512938)
         );
  XNOR2_X1 U106 ( .A(n445), .B(n466), .ZN(SUM[29]) );
  AND2_X1 U107 ( .A1(n364), .A2(n360), .ZN(n466) );
  NAND2_X1 U108 ( .A1(n326), .A2(n335), .ZN(n347) );
  NAND2_X1 U109 ( .A1(n303), .A2(n305), .ZN(n322) );
  NAND2_X1 U110 ( .A1(n307), .A2(n306), .ZN(n325) );
  NAND2_X1 U111 ( .A1(n328), .A2(n337), .ZN(n342) );
  NAND2_X1 U112 ( .A1(n284), .A2(n282), .ZN(n295) );
  NAND2_X1 U113 ( .A1(net512908), .A2(net512907), .ZN(n388) );
  NAND2_X1 U114 ( .A1(n363), .A2(n359), .ZN(n381) );
  AND2_X1 U115 ( .A1(net512987), .A2(net513003), .ZN(n19) );
  NAND2_X1 U116 ( .A1(net512905), .A2(net512901), .ZN(n384) );
  NAND2_X1 U117 ( .A1(n117), .A2(n116), .ZN(n18) );
  OAI21_X1 U118 ( .B1(n165), .B2(n548), .A(n449), .ZN(n164) );
  INV_X1 U119 ( .A(n307), .ZN(n517) );
  INV_X1 U120 ( .A(net512870), .ZN(n542) );
  AOI21_X1 U121 ( .B1(n402), .B2(net512987), .A(n543), .ZN(n401) );
  INV_X1 U122 ( .A(net512866), .ZN(n505) );
  OAI21_X1 U123 ( .B1(n476), .B2(n529), .A(n188), .ZN(n198) );
  INV_X1 U124 ( .A(n202), .ZN(n476) );
  OAI21_X1 U125 ( .B1(n475), .B2(n525), .A(n214), .ZN(n224) );
  INV_X1 U126 ( .A(n228), .ZN(n475) );
  OAI21_X1 U127 ( .B1(n478), .B2(n533), .A(n156), .ZN(n172) );
  INV_X1 U128 ( .A(n176), .ZN(n478) );
  OAI21_X1 U129 ( .B1(n477), .B2(n538), .A(n135), .ZN(n144) );
  AOI21_X1 U130 ( .B1(n423), .B2(n424), .A(n425), .ZN(n94) );
  OAI21_X1 U131 ( .B1(n207), .B2(n481), .A(n209), .ZN(n205) );
  NAND4_X1 U132 ( .A1(n219), .A2(n220), .A3(n218), .A4(n221), .ZN(n207) );
  AOI21_X1 U133 ( .B1(n210), .B2(n211), .A(n73), .ZN(n209) );
  OAI211_X1 U134 ( .C1(n525), .C2(n213), .A(n214), .B(n215), .ZN(n211) );
  OAI21_X1 U135 ( .B1(n540), .B2(n480), .A(n187), .ZN(n202) );
  INV_X1 U136 ( .A(n193), .ZN(n540) );
  OAI21_X1 U137 ( .B1(n541), .B2(n481), .A(n213), .ZN(n228) );
  INV_X1 U138 ( .A(n219), .ZN(n541) );
  OAI21_X1 U139 ( .B1(n181), .B2(n480), .A(n183), .ZN(n179) );
  NAND4_X1 U140 ( .A1(n193), .A2(n194), .A3(n192), .A4(n195), .ZN(n181) );
  AOI21_X1 U141 ( .B1(n184), .B2(n185), .A(n74), .ZN(n183) );
  OAI211_X1 U142 ( .C1(n529), .C2(n187), .A(n188), .B(n189), .ZN(n185) );
  OAI21_X1 U143 ( .B1(n539), .B2(n479), .A(n155), .ZN(n176) );
  INV_X1 U144 ( .A(n161), .ZN(n539) );
  OAI21_X1 U145 ( .B1(n149), .B2(n479), .A(n151), .ZN(n147) );
  NAND4_X1 U146 ( .A1(n161), .A2(n162), .A3(n160), .A4(n163), .ZN(n149) );
  AOI21_X1 U147 ( .B1(n152), .B2(n153), .A(n75), .ZN(n151) );
  OAI211_X1 U148 ( .C1(n533), .C2(n155), .A(n156), .B(n157), .ZN(n153) );
  OAI211_X1 U149 ( .C1(net537302), .C2(net513003), .A(net513004), .B(net513005), .ZN(n39) );
  NOR2_X1 U150 ( .A1(n513), .A2(n514), .ZN(n366) );
  INV_X1 U151 ( .A(n354), .ZN(n514) );
  NAND2_X1 U152 ( .A1(n276), .A2(n275), .ZN(n285) );
  OAI211_X1 U153 ( .C1(n516), .C2(n335), .A(n336), .B(n337), .ZN(n333) );
  NOR2_X1 U154 ( .A1(n504), .A2(n503), .ZN(n383) );
  XNOR2_X1 U155 ( .A(n450), .B(n229), .ZN(SUM[4]) );
  OAI21_X1 U156 ( .B1(n12), .B2(n274), .A(n275), .ZN(n251) );
  AND3_X1 U157 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n12) );
  NAND2_X1 U158 ( .A1(n276), .A2(n277), .ZN(n274) );
  NAND2_X1 U160 ( .A1(n281), .A2(n282), .ZN(n279) );
  NAND4_X1 U161 ( .A1(net512908), .A2(net512903), .A3(net512905), .A4(
        net512899), .ZN(net512810) );
  NAND4_X1 U162 ( .A1(net512943), .A2(net512944), .A3(net512936), .A4(
        net512937), .ZN(net512808) );
  NOR2_X1 U163 ( .A1(n508), .A2(n507), .ZN(net512876) );
  INV_X1 U164 ( .A(net512863), .ZN(n508) );
  AND3_X1 U165 ( .A1(net512905), .A2(n32), .A3(net512903), .ZN(n9) );
  NAND2_X1 U166 ( .A1(net512906), .A2(net512907), .ZN(n32) );
  XNOR2_X1 U167 ( .A(n234), .B(n233), .ZN(SUM[48]) );
  NAND2_X1 U168 ( .A1(n219), .A2(n213), .ZN(n234) );
  XNOR2_X1 U169 ( .A(n293), .B(n292), .ZN(SUM[41]) );
  NAND2_X1 U170 ( .A1(n278), .A2(n281), .ZN(n293) );
  XNOR2_X1 U171 ( .A(n345), .B(n344), .ZN(SUM[33]) );
  XNOR2_X1 U172 ( .A(n203), .B(n202), .ZN(SUM[53]) );
  NAND2_X1 U173 ( .A1(n194), .A2(n188), .ZN(n203) );
  XNOR2_X1 U174 ( .A(n206), .B(n205), .ZN(SUM[52]) );
  NAND2_X1 U175 ( .A1(n193), .A2(n187), .ZN(n206) );
  XNOR2_X1 U176 ( .A(n200), .B(n198), .ZN(SUM[54]) );
  NAND2_X1 U177 ( .A1(n192), .A2(n189), .ZN(n200) );
  XNOR2_X1 U178 ( .A(n231), .B(n228), .ZN(SUM[49]) );
  NAND2_X1 U179 ( .A1(n220), .A2(n214), .ZN(n231) );
  XNOR2_X1 U180 ( .A(n226), .B(n224), .ZN(SUM[50]) );
  NAND2_X1 U181 ( .A1(n218), .A2(n215), .ZN(n226) );
  XNOR2_X1 U182 ( .A(n272), .B(n271), .ZN(SUM[44]) );
  NAND2_X1 U183 ( .A1(n259), .A2(n246), .ZN(n272) );
  XNOR2_X1 U184 ( .A(n289), .B(n288), .ZN(SUM[42]) );
  NAND2_X1 U185 ( .A1(n280), .A2(n277), .ZN(n289) );
  XNOR2_X1 U186 ( .A(n266), .B(n265), .ZN(SUM[46]) );
  NAND2_X1 U187 ( .A1(n243), .A2(n247), .ZN(n266) );
  XNOR2_X1 U188 ( .A(n180), .B(n179), .ZN(SUM[56]) );
  NAND2_X1 U189 ( .A1(n161), .A2(n155), .ZN(n180) );
  XNOR2_X1 U190 ( .A(n177), .B(n176), .ZN(SUM[57]) );
  NAND2_X1 U191 ( .A1(n162), .A2(n156), .ZN(n177) );
  XNOR2_X1 U192 ( .A(n174), .B(n172), .ZN(SUM[58]) );
  NAND2_X1 U193 ( .A1(n160), .A2(n157), .ZN(n174) );
  XNOR2_X1 U194 ( .A(n145), .B(n144), .ZN(SUM[61]) );
  NAND2_X1 U195 ( .A1(n136), .A2(n134), .ZN(n145) );
  XNOR2_X1 U196 ( .A(n269), .B(n268), .ZN(SUM[45]) );
  NAND2_X1 U197 ( .A1(n260), .A2(n248), .ZN(n269) );
  XNOR2_X1 U198 ( .A(n148), .B(n147), .ZN(SUM[60]) );
  NAND2_X1 U199 ( .A1(n146), .A2(n135), .ZN(n148) );
  XNOR2_X1 U200 ( .A(n142), .B(n141), .ZN(SUM[62]) );
  NAND2_X1 U201 ( .A1(n137), .A2(n131), .ZN(n142) );
  XNOR2_X1 U202 ( .A(n138), .B(n139), .ZN(SUM[63]) );
  NAND2_X1 U203 ( .A1(n130), .A2(n126), .ZN(n139) );
  NAND2_X1 U204 ( .A1(n131), .A2(n140), .ZN(n138) );
  NAND2_X1 U205 ( .A1(n141), .A2(n137), .ZN(n140) );
  XNOR2_X1 U206 ( .A(n222), .B(n223), .ZN(SUM[51]) );
  NOR2_X1 U207 ( .A1(n528), .A2(n73), .ZN(n223) );
  AOI21_X1 U208 ( .B1(n218), .B2(n224), .A(n527), .ZN(n222) );
  INV_X1 U209 ( .A(n215), .ZN(n527) );
  XNOR2_X1 U210 ( .A(net537536), .B(net512961), .ZN(SUM[17]) );
  NAND2_X1 U211 ( .A1(net512944), .A2(n43), .ZN(net512961) );
  OAI211_X1 U212 ( .C1(net512962), .C2(n448), .A(net512964), .B(n42), .ZN(
        net537536) );
  AOI21_X1 U213 ( .B1(n39), .B2(n38), .A(n494), .ZN(n21) );
  NAND2_X1 U214 ( .A1(net512936), .A2(net512942), .ZN(net512956) );
  OAI21_X1 U215 ( .B1(n400), .B2(n489), .A(n47), .ZN(net538396) );
  AOI21_X1 U216 ( .B1(n402), .B2(net512987), .A(n543), .ZN(n47) );
  OAI211_X1 U217 ( .C1(n523), .C2(n246), .A(n247), .B(n248), .ZN(n239) );
  XNOR2_X1 U218 ( .A(n196), .B(n197), .ZN(SUM[55]) );
  NOR2_X1 U219 ( .A1(n532), .A2(n74), .ZN(n197) );
  AOI21_X1 U220 ( .B1(n192), .B2(n198), .A(n531), .ZN(n196) );
  INV_X1 U221 ( .A(n189), .ZN(n531) );
  XNOR2_X1 U222 ( .A(n170), .B(n171), .ZN(SUM[59]) );
  NOR2_X1 U223 ( .A1(n536), .A2(n75), .ZN(n171) );
  AOI21_X1 U224 ( .B1(n160), .B2(n172), .A(n535), .ZN(n170) );
  INV_X1 U225 ( .A(n157), .ZN(n535) );
  XNOR2_X1 U226 ( .A(n314), .B(n315), .ZN(SUM[39]) );
  OAI21_X1 U227 ( .B1(n98), .B2(n99), .A(n100), .ZN(n97) );
  NAND2_X1 U228 ( .A1(n101), .A2(n102), .ZN(n99) );
  XNOR2_X1 U229 ( .A(n262), .B(n263), .ZN(SUM[47]) );
  NAND2_X1 U230 ( .A1(n242), .A2(n244), .ZN(n262) );
  NAND2_X1 U231 ( .A1(n264), .A2(n247), .ZN(n263) );
  NAND2_X1 U232 ( .A1(n243), .A2(n265), .ZN(n264) );
  AND2_X1 U233 ( .A1(n411), .A2(n407), .ZN(n53) );
  OR2_X1 U234 ( .A1(net512990), .A2(n497), .ZN(net512964) );
  INV_X1 U235 ( .A(net512943), .ZN(n497) );
  AOI21_X1 U236 ( .B1(n38), .B2(n39), .A(n494), .ZN(net512990) );
  NAND2_X1 U237 ( .A1(n116), .A2(n449), .ZN(n103) );
  NAND4_X1 U238 ( .A1(n284), .A2(n278), .A3(n280), .A4(n275), .ZN(n254) );
  XNOR2_X1 U239 ( .A(n395), .B(n396), .ZN(SUM[15]) );
  NAND2_X1 U240 ( .A1(net513001), .A2(net512986), .ZN(n396) );
  NAND2_X1 U241 ( .A1(n493), .A2(net512989), .ZN(n397) );
  AND2_X1 U242 ( .A1(net512903), .A2(net512906), .ZN(n467) );
  NOR2_X1 U243 ( .A1(n528), .A2(n526), .ZN(n210) );
  INV_X1 U244 ( .A(n218), .ZN(n526) );
  NOR2_X1 U245 ( .A1(n532), .A2(n530), .ZN(n184) );
  INV_X1 U246 ( .A(n192), .ZN(n530) );
  NOR2_X1 U247 ( .A1(n536), .A2(n534), .ZN(n152) );
  INV_X1 U248 ( .A(n160), .ZN(n534) );
  NAND2_X1 U249 ( .A1(n270), .A2(n246), .ZN(n268) );
  NAND2_X1 U250 ( .A1(n271), .A2(n259), .ZN(n270) );
  NOR2_X1 U251 ( .A1(n105), .A2(n548), .ZN(n98) );
  NAND2_X1 U252 ( .A1(n107), .A2(n108), .ZN(n105) );
  INV_X1 U253 ( .A(net537302), .ZN(n492) );
  NAND2_X1 U254 ( .A1(n143), .A2(n134), .ZN(n141) );
  NAND2_X1 U255 ( .A1(n136), .A2(n144), .ZN(n143) );
  INV_X1 U256 ( .A(n106), .ZN(n548) );
  OAI21_X1 U257 ( .B1(n103), .B2(n106), .A(n104), .ZN(n114) );
  NAND2_X1 U258 ( .A1(n374), .A2(n390), .ZN(n168) );
  AND2_X1 U259 ( .A1(n427), .A2(n411), .ZN(n67) );
  NAND2_X1 U260 ( .A1(net512943), .A2(n25), .ZN(net512962) );
  NAND2_X1 U261 ( .A1(n115), .A2(n116), .ZN(n104) );
  OAI211_X1 U262 ( .C1(net538262), .C2(net512962), .A(net512964), .B(n42), 
        .ZN(net512958) );
  INV_X1 U263 ( .A(n110), .ZN(n490) );
  AND4_X1 U264 ( .A1(n492), .A2(net512986), .A3(net512987), .A4(net512989), 
        .ZN(n25) );
  AND2_X1 U265 ( .A1(n427), .A2(n411), .ZN(n64) );
  NAND2_X1 U266 ( .A1(net512987), .A2(n59), .ZN(n400) );
  AND4_X1 U267 ( .A1(n326), .A2(n327), .A3(n328), .A4(n329), .ZN(n71) );
  INV_X1 U268 ( .A(net513001), .ZN(n494) );
  INV_X1 U269 ( .A(net512944), .ZN(n498) );
  INV_X1 U270 ( .A(n221), .ZN(n528) );
  INV_X1 U271 ( .A(n195), .ZN(n532) );
  INV_X1 U272 ( .A(n163), .ZN(n536) );
  INV_X1 U273 ( .A(n146), .ZN(n538) );
  INV_X1 U274 ( .A(n220), .ZN(n525) );
  INV_X1 U275 ( .A(n194), .ZN(n529) );
  INV_X1 U276 ( .A(n162), .ZN(n533) );
  INV_X1 U277 ( .A(n260), .ZN(n523) );
  INV_X1 U278 ( .A(net513003), .ZN(n543) );
  AND4_X1 U279 ( .A1(n259), .A2(n260), .A3(n243), .A4(n244), .ZN(n72) );
  AND2_X1 U280 ( .A1(n100), .A2(n117), .ZN(n423) );
  AND2_X1 U281 ( .A1(n305), .A2(n306), .ZN(n11) );
  OAI21_X1 U282 ( .B1(n548), .B2(n87), .A(n439), .ZN(n85) );
  NOR2_X1 U283 ( .A1(n51), .A2(n490), .ZN(n84) );
  INV_X1 U284 ( .A(net513004), .ZN(n493) );
  XNOR2_X1 U285 ( .A(n468), .B(n469), .ZN(SUM[6]) );
  NAND2_X1 U286 ( .A1(n111), .A2(n112), .ZN(n468) );
  NAND2_X1 U287 ( .A1(n102), .A2(n100), .ZN(n469) );
  INV_X1 U288 ( .A(n303), .ZN(n519) );
  OAI21_X1 U289 ( .B1(n485), .B2(n521), .A(n281), .ZN(n288) );
  INV_X1 U290 ( .A(n278), .ZN(n521) );
  INV_X1 U291 ( .A(n292), .ZN(n485) );
  INV_X1 U292 ( .A(net512903), .ZN(n500) );
  AND2_X1 U293 ( .A1(n243), .A2(n244), .ZN(n240) );
  NAND2_X1 U294 ( .A1(n64), .A2(n426), .ZN(n415) );
  NAND2_X1 U295 ( .A1(n428), .A2(n110), .ZN(n426) );
  INV_X1 U296 ( .A(n411), .ZN(n545) );
  INV_X1 U297 ( .A(net512899), .ZN(n503) );
  NAND2_X1 U298 ( .A1(n547), .A2(n491), .ZN(n111) );
  INV_X1 U299 ( .A(net512862), .ZN(n507) );
  INV_X1 U300 ( .A(n356), .ZN(n513) );
  OAI21_X1 U301 ( .B1(n484), .B2(n523), .A(n248), .ZN(n265) );
  INV_X1 U302 ( .A(n268), .ZN(n484) );
  INV_X1 U303 ( .A(n242), .ZN(n524) );
  INV_X1 U304 ( .A(net512864), .ZN(n506) );
  INV_X1 U305 ( .A(net512901), .ZN(n502) );
  INV_X1 U306 ( .A(n361), .ZN(n512) );
  INV_X1 U307 ( .A(n428), .ZN(n546) );
  XNOR2_X1 U308 ( .A(n372), .B(n313), .ZN(SUM[2]) );
  NAND2_X1 U309 ( .A1(n377), .A2(n312), .ZN(n372) );
  XNOR2_X1 U310 ( .A(n308), .B(n309), .ZN(SUM[3]) );
  OAI21_X1 U311 ( .B1(n551), .B2(n549), .A(n312), .ZN(n309) );
  INV_X1 U312 ( .A(n377), .ZN(n549) );
  XNOR2_X1 U313 ( .A(n389), .B(n553), .ZN(SUM[1]) );
  NAND2_X1 U314 ( .A1(n375), .A2(n374), .ZN(n389) );
  NAND2_X1 U315 ( .A1(n555), .A2(n550), .ZN(n377) );
  NAND2_X1 U316 ( .A1(n554), .A2(n552), .ZN(n375) );
  AOI21_X1 U317 ( .B1(n127), .B2(n128), .A(n129), .ZN(n124) );
  AND2_X1 U318 ( .A1(n136), .A2(n137), .ZN(n127) );
  NAND2_X1 U319 ( .A1(n130), .A2(n131), .ZN(n129) );
  OAI211_X1 U320 ( .C1(n477), .C2(n538), .A(n134), .B(n135), .ZN(n128) );
  NAND2_X1 U321 ( .A1(n554), .A2(n552), .ZN(n91) );
  NAND2_X1 U322 ( .A1(n373), .A2(n374), .ZN(n313) );
  NAND2_X1 U323 ( .A1(n375), .A2(n553), .ZN(n373) );
  NAND2_X1 U324 ( .A1(n374), .A2(n390), .ZN(n92) );
  INV_X1 U325 ( .A(n390), .ZN(n553) );
  NAND2_X1 U326 ( .A1(n555), .A2(n550), .ZN(n167) );
  INV_X1 U327 ( .A(n126), .ZN(n537) );
  AND3_X1 U328 ( .A1(B[8]), .A2(n411), .A3(A[8]), .ZN(n405) );
  NOR2_X1 U329 ( .A1(B[13]), .A2(A[13]), .ZN(net537302) );
  OR2_X1 U330 ( .A1(B[12]), .A2(A[12]), .ZN(net512987) );
  NAND2_X1 U331 ( .A1(B[3]), .A2(A[3]), .ZN(n106) );
  NAND2_X1 U332 ( .A1(n391), .A2(n407), .ZN(n413) );
  NAND2_X1 U333 ( .A1(B[7]), .A2(A[7]), .ZN(n110) );
  OR2_X1 U334 ( .A1(B[50]), .A2(A[50]), .ZN(n218) );
  OR2_X1 U335 ( .A1(B[54]), .A2(A[54]), .ZN(n192) );
  OR2_X1 U336 ( .A1(B[58]), .A2(A[58]), .ZN(n160) );
  NAND2_X1 U337 ( .A1(B[13]), .A2(A[13]), .ZN(net513004) );
  NAND2_X1 U338 ( .A1(B[46]), .A2(A[46]), .ZN(n247) );
  NAND2_X1 U339 ( .A1(B[44]), .A2(A[44]), .ZN(n246) );
  NAND2_X1 U340 ( .A1(B[61]), .A2(A[61]), .ZN(n134) );
  NAND2_X1 U341 ( .A1(B[20]), .A2(A[20]), .ZN(net512907) );
  NAND2_X1 U342 ( .A1(B[18]), .A2(A[18]), .ZN(net512942) );
  NAND2_X1 U343 ( .A1(B[53]), .A2(A[53]), .ZN(n188) );
  NAND2_X1 U344 ( .A1(B[49]), .A2(A[49]), .ZN(n214) );
  NAND2_X1 U345 ( .A1(B[50]), .A2(A[50]), .ZN(n215) );
  NAND2_X1 U346 ( .A1(B[52]), .A2(A[52]), .ZN(n187) );
  NAND2_X1 U347 ( .A1(B[48]), .A2(A[48]), .ZN(n213) );
  NAND2_X1 U348 ( .A1(B[45]), .A2(A[45]), .ZN(n248) );
  NAND2_X1 U349 ( .A1(B[57]), .A2(A[57]), .ZN(n156) );
  NAND2_X1 U350 ( .A1(B[62]), .A2(A[62]), .ZN(n131) );
  NAND2_X1 U351 ( .A1(B[54]), .A2(A[54]), .ZN(n189) );
  NAND2_X1 U352 ( .A1(B[58]), .A2(A[58]), .ZN(n157) );
  NAND2_X1 U353 ( .A1(B[56]), .A2(A[56]), .ZN(n155) );
  NAND2_X1 U354 ( .A1(B[8]), .A2(A[8]), .ZN(n428) );
  NAND2_X1 U355 ( .A1(B[60]), .A2(A[60]), .ZN(n135) );
  NAND2_X1 U356 ( .A1(B[41]), .A2(A[41]), .ZN(n281) );
  NAND2_X1 U357 ( .A1(B[22]), .A2(A[22]), .ZN(net512901) );
  NAND2_X1 U358 ( .A1(B[30]), .A2(A[30]), .ZN(n361) );
  OR2_X1 U359 ( .A1(B[46]), .A2(A[46]), .ZN(n243) );
  OR2_X1 U360 ( .A1(B[21]), .A2(A[21]), .ZN(net512903) );
  OR2_X1 U361 ( .A1(B[41]), .A2(A[41]), .ZN(n278) );
  NAND2_X1 U362 ( .A1(B[40]), .A2(A[40]), .ZN(n282) );
  NAND2_X1 U363 ( .A1(B[42]), .A2(A[42]), .ZN(n277) );
  NAND2_X1 U364 ( .A1(A[5]), .A2(B[5]), .ZN(n117) );
  NAND2_X1 U365 ( .A1(B[32]), .A2(A[32]), .ZN(n335) );
  NAND2_X1 U366 ( .A1(B[34]), .A2(A[34]), .ZN(n337) );
  NAND2_X1 U367 ( .A1(B[24]), .A2(A[24]), .ZN(net512870) );
  NAND2_X1 U368 ( .A1(B[12]), .A2(A[12]), .ZN(net513003) );
  NAND2_X1 U369 ( .A1(B[21]), .A2(A[21]), .ZN(net512906) );
  OR2_X1 U370 ( .A1(B[22]), .A2(A[22]), .ZN(net512905) );
  OR2_X1 U371 ( .A1(B[43]), .A2(A[43]), .ZN(n275) );
  NAND2_X1 U372 ( .A1(B[33]), .A2(A[33]), .ZN(n336) );
  NAND2_X1 U373 ( .A1(B[11]), .A2(n433), .ZN(n391) );
  OR2_X1 U374 ( .A1(B[42]), .A2(A[42]), .ZN(n280) );
  OR2_X1 U375 ( .A1(B[18]), .A2(A[18]), .ZN(net512936) );
  OR2_X1 U376 ( .A1(B[23]), .A2(A[23]), .ZN(net512899) );
  NAND2_X1 U377 ( .A1(B[9]), .A2(A[9]), .ZN(n80) );
  OR2_X1 U378 ( .A1(B[37]), .A2(A[37]), .ZN(n303) );
  NAND2_X1 U379 ( .A1(B[36]), .A2(A[36]), .ZN(n306) );
  NAND2_X1 U380 ( .A1(B[38]), .A2(A[38]), .ZN(n301) );
  NAND2_X1 U381 ( .A1(B[37]), .A2(A[37]), .ZN(n305) );
  NAND2_X1 U382 ( .A1(B[28]), .A2(A[28]), .ZN(n359) );
  NAND2_X1 U383 ( .A1(B[14]), .A2(A[14]), .ZN(net513005) );
  NAND2_X1 U384 ( .A1(B[6]), .A2(A[6]), .ZN(n100) );
  OR2_X1 U385 ( .A1(B[49]), .A2(A[49]), .ZN(n220) );
  OR2_X1 U386 ( .A1(B[53]), .A2(A[53]), .ZN(n194) );
  OR2_X1 U387 ( .A1(B[57]), .A2(A[57]), .ZN(n162) );
  OR2_X1 U388 ( .A1(B[45]), .A2(A[45]), .ZN(n260) );
  OR2_X1 U389 ( .A1(B[44]), .A2(A[44]), .ZN(n259) );
  OR2_X1 U390 ( .A1(B[52]), .A2(A[52]), .ZN(n193) );
  OR2_X1 U391 ( .A1(B[48]), .A2(A[48]), .ZN(n219) );
  OR2_X1 U392 ( .A1(B[56]), .A2(A[56]), .ZN(n161) );
  NAND2_X1 U393 ( .A1(B[47]), .A2(A[47]), .ZN(n242) );
  OR2_X1 U394 ( .A1(B[47]), .A2(A[47]), .ZN(n244) );
  OR2_X1 U395 ( .A1(B[19]), .A2(A[19]), .ZN(net512937) );
  NAND2_X1 U396 ( .A1(B[63]), .A2(A[63]), .ZN(n130) );
  NAND2_X1 U397 ( .A1(B[19]), .A2(A[19]), .ZN(net512935) );
  OR2_X1 U398 ( .A1(B[34]), .A2(A[34]), .ZN(n328) );
  OR2_X1 U399 ( .A1(B[62]), .A2(A[62]), .ZN(n137) );
  NAND2_X1 U400 ( .A1(B[25]), .A2(A[25]), .ZN(net512869) );
  OR2_X1 U401 ( .A1(B[25]), .A2(A[25]), .ZN(net512866) );
  OR2_X1 U402 ( .A1(B[36]), .A2(A[36]), .ZN(n307) );
  OR2_X1 U403 ( .A1(B[61]), .A2(A[61]), .ZN(n136) );
  OR2_X1 U404 ( .A1(B[20]), .A2(A[20]), .ZN(net512908) );
  OR2_X1 U405 ( .A1(B[40]), .A2(A[40]), .ZN(n284) );
  NAND2_X1 U406 ( .A1(B[23]), .A2(A[23]), .ZN(net512900) );
  OR2_X1 U407 ( .A1(B[38]), .A2(A[38]), .ZN(n304) );
  AND2_X1 U408 ( .A1(B[51]), .A2(A[51]), .ZN(n73) );
  AND2_X1 U409 ( .A1(B[55]), .A2(A[55]), .ZN(n74) );
  AND2_X1 U410 ( .A1(B[59]), .A2(A[59]), .ZN(n75) );
  OR2_X1 U411 ( .A1(B[27]), .A2(A[27]), .ZN(net512862) );
  OR2_X1 U412 ( .A1(B[31]), .A2(A[31]), .ZN(n356) );
  OR2_X1 U413 ( .A1(B[51]), .A2(A[51]), .ZN(n221) );
  OR2_X1 U414 ( .A1(B[55]), .A2(A[55]), .ZN(n195) );
  OR2_X1 U415 ( .A1(B[59]), .A2(A[59]), .ZN(n163) );
  OR2_X1 U416 ( .A1(B[32]), .A2(A[32]), .ZN(n326) );
  OR2_X1 U417 ( .A1(B[24]), .A2(A[24]), .ZN(net512871) );
  OR2_X1 U418 ( .A1(B[28]), .A2(A[28]), .ZN(n363) );
  OR2_X1 U419 ( .A1(B[63]), .A2(A[63]), .ZN(n126) );
  OR2_X1 U420 ( .A1(B[60]), .A2(A[60]), .ZN(n146) );
  OR2_X1 U421 ( .A1(A[8]), .A2(B[8]), .ZN(n82) );
  OR2_X1 U422 ( .A1(B[35]), .A2(A[35]), .ZN(n329) );
  OR2_X1 U423 ( .A1(B[33]), .A2(A[33]), .ZN(n327) );
  OR2_X1 U424 ( .A1(B[8]), .A2(A[8]), .ZN(n427) );
  OR2_X1 U425 ( .A1(B[7]), .A2(A[7]), .ZN(n3) );
  OR2_X1 U426 ( .A1(B[15]), .A2(A[15]), .ZN(n41) );
  NAND2_X1 U427 ( .A1(B[2]), .A2(n437), .ZN(n312) );
  INV_X1 U428 ( .A(n437), .ZN(n550) );
  INV_X1 U429 ( .A(B[2]), .ZN(n555) );
  INV_X1 U430 ( .A(A[1]), .ZN(n552) );
  OR2_X1 U431 ( .A1(B[0]), .A2(A[0]), .ZN(n429) );
  NAND2_X1 U432 ( .A1(B[1]), .A2(A[1]), .ZN(n374) );
  NAND2_X1 U433 ( .A1(B[0]), .A2(A[0]), .ZN(n390) );
  INV_X1 U434 ( .A(B[1]), .ZN(n554) );
  NAND2_X1 U435 ( .A1(n59), .A2(n95), .ZN(n403) );
  INV_X1 U436 ( .A(n95), .ZN(n489) );
  OAI21_X1 U437 ( .B1(n489), .B2(n400), .A(n401), .ZN(n398) );
  XNOR2_X1 U438 ( .A(n17), .B(n18), .ZN(SUM[5]) );
  NAND2_X1 U439 ( .A1(B[27]), .A2(A[27]), .ZN(net512863) );
  NAND2_X1 U440 ( .A1(net512866), .A2(net512869), .ZN(net512889) );
  NAND2_X1 U441 ( .A1(net512869), .A2(net512870), .ZN(net512867) );
  AND2_X1 U442 ( .A1(n60), .A2(n408), .ZN(n56) );
  NAND2_X1 U443 ( .A1(n80), .A2(n408), .ZN(n406) );
  NAND2_X1 U444 ( .A1(B[26]), .A2(A[26]), .ZN(net512864) );
  NAND2_X1 U445 ( .A1(B[16]), .A2(A[16]), .ZN(n42) );
  CLKBUF_X1 U446 ( .A(n283), .Z(n470) );
  OAI21_X1 U447 ( .B1(n483), .B2(n519), .A(n305), .ZN(n317) );
  XNOR2_X1 U448 ( .A(n295), .B(n470), .ZN(SUM[40]) );
  NAND2_X1 U449 ( .A1(n522), .A2(n470), .ZN(n273) );
  OAI21_X1 U450 ( .B1(n486), .B2(n261), .A(n252), .ZN(n283) );
  OAI21_X1 U451 ( .B1(n517), .B2(n486), .A(n306), .ZN(n321) );
  XNOR2_X1 U452 ( .A(n473), .B(net512889), .ZN(SUM[25]) );
  AND2_X1 U453 ( .A1(n167), .A2(n438), .ZN(n8) );
  NAND4_X1 U454 ( .A1(n91), .A2(n167), .A3(n168), .A4(n438), .ZN(n166) );
  NAND2_X1 U455 ( .A1(n438), .A2(n106), .ZN(n308) );
  NOR2_X1 U456 ( .A1(B[10]), .A2(A[10]), .ZN(n44) );
  OR2_X1 U457 ( .A1(B[10]), .A2(A[10]), .ZN(n60) );
  NAND2_X1 U458 ( .A1(A[10]), .A2(B[10]), .ZN(n408) );
  INV_X1 U459 ( .A(n324), .ZN(n486) );
  XNOR2_X1 U460 ( .A(n325), .B(n324), .ZN(SUM[36]) );
  NAND4_X1 U461 ( .A1(n518), .A2(n522), .A3(n71), .A4(n72), .ZN(n235) );
  XNOR2_X1 U462 ( .A(net537535), .B(net512956), .ZN(SUM[18]) );
  NAND2_X1 U463 ( .A1(B[29]), .A2(A[29]), .ZN(n360) );
  OR2_X1 U464 ( .A1(B[29]), .A2(A[29]), .ZN(n364) );
  NAND2_X1 U465 ( .A1(B[17]), .A2(A[17]), .ZN(n43) );
  OAI21_X1 U466 ( .B1(n444), .B2(n442), .A(n412), .ZN(n58) );
  OAI21_X1 U467 ( .B1(n45), .B2(n442), .A(n412), .ZN(n95) );
  NAND2_X1 U468 ( .A1(n301), .A2(n316), .ZN(n315) );
  XNOR2_X1 U469 ( .A(n285), .B(n286), .ZN(SUM[43]) );
  NAND2_X1 U470 ( .A1(B[43]), .A2(A[43]), .ZN(n276) );
  NAND2_X1 U471 ( .A1(net512953), .A2(net512936), .ZN(n23) );
  NAND2_X1 U472 ( .A1(n277), .A2(n287), .ZN(n286) );
  OAI21_X1 U473 ( .B1(n297), .B2(n298), .A(n299), .ZN(n252) );
  NAND2_X1 U474 ( .A1(n449), .A2(n118), .ZN(n229) );
  NAND2_X1 U475 ( .A1(n118), .A2(n117), .ZN(n115) );
  NAND2_X1 U476 ( .A1(net512868), .A2(net512864), .ZN(net512883) );
  AND3_X1 U477 ( .A1(net512866), .A2(net512867), .A3(net512868), .ZN(n10) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(SUM[11]) );
  OAI21_X1 U479 ( .B1(n68), .B2(n44), .A(n408), .ZN(n414) );
  OAI211_X1 U480 ( .C1(n405), .C2(n406), .A(n60), .B(n407), .ZN(n392) );
  OAI21_X1 U481 ( .B1(n445), .B2(n510), .A(n360), .ZN(n52) );
  OAI21_X1 U482 ( .B1(n54), .B2(n510), .A(n360), .ZN(n369) );
  OAI211_X1 U483 ( .C1(n510), .C2(n359), .A(n360), .B(n361), .ZN(n357) );
  INV_X1 U484 ( .A(n364), .ZN(n510) );
  OR2_X1 U485 ( .A1(B[7]), .A2(A[7]), .ZN(n109) );
  XNOR2_X1 U486 ( .A(n76), .B(n77), .ZN(SUM[9]) );
  AOI21_X1 U487 ( .B1(n81), .B2(n82), .A(n546), .ZN(n76) );
  NAND2_X1 U488 ( .A1(n356), .A2(n355), .ZN(n353) );
  INV_X1 U489 ( .A(net512900), .ZN(n504) );
  NAND2_X1 U490 ( .A1(net512900), .A2(net512901), .ZN(n31) );
  NAND2_X1 U491 ( .A1(n327), .A2(n336), .ZN(n345) );
  INV_X1 U492 ( .A(n327), .ZN(n516) );
  AOI21_X1 U493 ( .B1(n423), .B2(n424), .A(n425), .ZN(n51) );
  NAND2_X1 U494 ( .A1(n3), .A2(n102), .ZN(n425) );
  AND2_X1 U495 ( .A1(n108), .A2(n62), .ZN(n45) );
  NOR2_X1 U496 ( .A1(n94), .A2(n490), .ZN(n412) );
  NAND2_X1 U497 ( .A1(n518), .A2(n256), .ZN(n253) );
  XNOR2_X1 U498 ( .A(n382), .B(n383), .ZN(SUM[23]) );
  OAI21_X1 U499 ( .B1(n496), .B2(net512934), .A(net512935), .ZN(net512827) );
  INV_X1 U500 ( .A(net512938), .ZN(n496) );
  NAND2_X1 U501 ( .A1(net512936), .A2(net512937), .ZN(net512934) );
  OAI21_X1 U502 ( .B1(n4), .B2(n500), .A(net512906), .ZN(n16) );
  NOR2_X1 U503 ( .A1(n11), .A2(n302), .ZN(n297) );
  XNOR2_X1 U504 ( .A(net512875), .B(net512876), .ZN(SUM[27]) );
  NAND2_X1 U505 ( .A1(n329), .A2(n332), .ZN(n338) );
  OAI21_X1 U507 ( .B1(n471), .B2(n498), .A(n43), .ZN(net537535) );
  OAI21_X1 U508 ( .B1(n471), .B2(n498), .A(n43), .ZN(net512953) );
  AND2_X1 U509 ( .A1(n391), .A2(n392), .ZN(net512977) );
  NAND2_X1 U510 ( .A1(n391), .A2(n392), .ZN(n402) );
  AOI21_X1 U511 ( .B1(n252), .B2(n253), .A(n254), .ZN(n249) );
  INV_X1 U512 ( .A(n254), .ZN(n522) );
  OAI21_X1 U513 ( .B1(n515), .B2(n331), .A(n332), .ZN(n256) );
  NAND2_X1 U514 ( .A1(n328), .A2(n329), .ZN(n331) );
  INV_X1 U515 ( .A(n333), .ZN(n515) );
  NAND2_X1 U516 ( .A1(B[39]), .A2(A[39]), .ZN(n300) );
  OR2_X1 U517 ( .A1(B[39]), .A2(A[39]), .ZN(n299) );
  XNOR2_X1 U518 ( .A(net512881), .B(net512883), .ZN(SUM[26]) );
  AOI21_X1 U519 ( .B1(net512881), .B2(net512868), .A(n506), .ZN(net512875) );
  AOI21_X1 U520 ( .B1(n30), .B2(net512871), .A(n542), .ZN(net537046) );
  NOR2_X1 U521 ( .A1(n113), .A2(n114), .ZN(n112) );
  NAND2_X1 U522 ( .A1(A[4]), .A2(B[4]), .ZN(n118) );
  NAND2_X1 U523 ( .A1(n304), .A2(n301), .ZN(n318) );
  NAND4_X1 U524 ( .A1(n307), .A2(n303), .A3(n304), .A4(n299), .ZN(n261) );
  NAND2_X1 U525 ( .A1(n303), .A2(n304), .ZN(n302) );
  INV_X1 U526 ( .A(n357), .ZN(n509) );
  NAND2_X1 U527 ( .A1(n294), .A2(n282), .ZN(n292) );
  NAND2_X1 U528 ( .A1(n300), .A2(n299), .ZN(n314) );
  NAND2_X1 U529 ( .A1(n300), .A2(n301), .ZN(n298) );
  XNOR2_X1 U530 ( .A(n398), .B(net513018), .ZN(SUM[13]) );
  AOI21_X1 U531 ( .B1(n398), .B2(n492), .A(n493), .ZN(n29) );
  XNOR2_X1 U532 ( .A(n16), .B(n384), .ZN(SUM[22]) );
  AOI21_X1 U533 ( .B1(n16), .B2(net512905), .A(n502), .ZN(n382) );
  XNOR2_X1 U534 ( .A(net537976), .B(n388), .ZN(SUM[20]) );
  AND2_X1 U535 ( .A1(n387), .A2(net512907), .ZN(n4) );
  NAND2_X1 U536 ( .A1(net537976), .A2(net512908), .ZN(n387) );
  NAND2_X1 U537 ( .A1(B[35]), .A2(A[35]), .ZN(n332) );
  NAND2_X1 U538 ( .A1(n84), .A2(n85), .ZN(n81) );
  INV_X1 U539 ( .A(n454), .ZN(n547) );
  AND2_X1 U540 ( .A1(n104), .A2(n453), .ZN(n107) );
  NAND2_X1 U541 ( .A1(n166), .A2(n453), .ZN(n165) );
  NAND2_X1 U542 ( .A1(n89), .A2(n453), .ZN(n87) );
  AND2_X1 U543 ( .A1(n106), .A2(n90), .ZN(n62) );
  INV_X1 U544 ( .A(net512958), .ZN(n471) );
  OR2_X1 U545 ( .A1(B[15]), .A2(A[15]), .ZN(net512986) );
  NAND2_X1 U546 ( .A1(A[15]), .A2(B[15]), .ZN(net513001) );
  NAND2_X1 U547 ( .A1(n164), .A2(n118), .ZN(n17) );
  XNOR2_X1 U548 ( .A(n380), .B(n381), .ZN(SUM[28]) );
  OAI21_X1 U549 ( .B1(n362), .B2(net512809), .A(net512825), .ZN(n350) );
  NOR2_X1 U550 ( .A1(net512809), .A2(net512810), .ZN(net512804) );
  NAND2_X1 U551 ( .A1(n380), .A2(n363), .ZN(n379) );
  NOR2_X1 U552 ( .A1(net512807), .A2(net512808), .ZN(net512806) );
  XNOR2_X1 U553 ( .A(n321), .B(n322), .ZN(SUM[37]) );
  INV_X1 U554 ( .A(n321), .ZN(n483) );
  INV_X1 U555 ( .A(net512829), .ZN(n499) );
  INV_X1 U556 ( .A(n451), .ZN(n473) );
  OAI21_X1 U557 ( .B1(net537046), .B2(n505), .A(net512869), .ZN(net512881) );
  OAI21_X1 U558 ( .B1(n474), .B2(net512810), .A(net512829), .ZN(n30) );
  XNOR2_X1 U559 ( .A(n365), .B(n366), .ZN(SUM[31]) );
  AOI21_X1 U560 ( .B1(n369), .B2(n355), .A(n512), .ZN(n365) );
  OAI21_X1 U561 ( .B1(n10), .B2(net512861), .A(net512862), .ZN(net512825) );
  NAND2_X1 U563 ( .A1(net512863), .A2(net512864), .ZN(net512861) );
  OAI21_X1 U564 ( .B1(n472), .B2(net512809), .A(net512825), .ZN(n380) );
  NAND4_X1 U565 ( .A1(net512871), .A2(net512866), .A3(net512868), .A4(
        net512862), .ZN(net512809) );
  NAND2_X1 U566 ( .A1(n280), .A2(n288), .ZN(n287) );
  NAND2_X1 U567 ( .A1(n283), .A2(n284), .ZN(n294) );
  INV_X1 U568 ( .A(n257), .ZN(n482) );
  XNOR2_X1 U569 ( .A(n342), .B(n341), .ZN(SUM[34]) );
  NAND2_X1 U570 ( .A1(n328), .A2(n341), .ZN(n340) );
  XNOR2_X1 U571 ( .A(n347), .B(n257), .ZN(SUM[32]) );
  AND2_X1 U572 ( .A1(n71), .A2(n257), .ZN(n69) );
  NAND2_X1 U573 ( .A1(B[31]), .A2(A[31]), .ZN(n354) );
  XNOR2_X1 U574 ( .A(n317), .B(n318), .ZN(SUM[38]) );
  NAND2_X1 U578 ( .A1(n304), .A2(n317), .ZN(n316) );
  AOI21_X1 U579 ( .B1(n511), .B2(n350), .A(n351), .ZN(n348) );
  OAI21_X1 U580 ( .B1(n509), .B2(n353), .A(n354), .ZN(n351) );
  INV_X1 U581 ( .A(net512807), .ZN(n511) );
  NAND2_X1 U582 ( .A1(n348), .A2(n349), .ZN(n257) );
  XNOR2_X1 U584 ( .A(n339), .B(n338), .ZN(SUM[35]) );
  NAND2_X1 U585 ( .A1(n340), .A2(n337), .ZN(n339) );
  OAI21_X1 U586 ( .B1(n487), .B2(n516), .A(n336), .ZN(n341) );
  INV_X1 U588 ( .A(n344), .ZN(n487) );
endmodule


module RCA_NBIT64_0 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_0_DW01_add_9 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_14_DW01_add_6 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net507395, net507383, net507382, net507370, net507360, net507358,
         net507352, net507347, net507346, net507341, net507340, net507318,
         net507302, net507301, net507300, net507296, net507283, net507282,
         net507280, net507279, net507278, net507122, net535421, net537206,
         net537591, net537590, net537652, net538645, net507312, net507291,
         net507349, net507345, net507343, net507339, net507367, net507344,
         net507338, net507295, net507313, net537017, net507348, net507297,
         net537128, net507336, net507314, net507307, net507306, net507290,
         net507287, net507286, net507285, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n26, n27, n29, n31,
         n33, n34, n36, n39, n40, n41, n44, n45, n46, n47, n48, n52, n53, n55,
         n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n72, n73, n74, n75, n77, n78, n79, n80, n82, n83, n85, n86, n87, n88,
         n89, n90, n93, n94, n97, n98, n100, n101, n102, n104, n105, n106,
         n107, n108, n109, n110, n112, n113, n114, n116, n117, n118, n121,
         n122, n123, n124, n125, n126, n129, n130, n131, n132, n134, n136,
         n137, n139, n140, n141, n143, n144, n145, n147, n148, n149, n152,
         n153, n154, n155, n156, n157, n158, n162, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n178, n180, n181,
         n182, n183, n184, n185, n186, n187, n189, n190, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n204, n205, n207,
         n208, n209, n210, n211, n213, n214, n215, n216, n217, n219, n221,
         n222, n223, n224, n225, n226, n227, n228, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n247, n248, n249, n250, n251, n252, n253, n256, n257, n258,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n288, n290, n291, n292, n293, n294, n295, n297, n298, n299,
         n301, n302, n303, n304, n305, n306, n307, n310, n311, n312, n314,
         n315, n316, n317, n318, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n336, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n358, n359, n361, n362, n363, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n378, n380, n381, n382, n383, n385, n386, n387, n388, n389, n390,
         n391, n392, n394, n395, n396, n397, n398, n400, n401, n404, n405,
         n406, n407, n408, n409, n410, n411, n413, n414, n415, n416, n417,
         n418, n419, n422, n423, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n436, n437, n439, n440, n441, n442, n443, n444,
         n447, n448, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568;

  AND2_X2 U4 ( .A1(B[4]), .A2(A[4]), .ZN(n46) );
  NAND3_X1 U71 ( .A1(net535421), .A2(net537017), .A3(n16), .ZN(net507278) );
  NAND3_X1 U114 ( .A1(n323), .A2(n461), .A3(n17), .ZN(net507301) );
  OR2_X2 U129 ( .A1(A[5]), .A2(B[5]), .ZN(n80) );
  OR2_X2 U319 ( .A1(A[7]), .A2(B[7]), .ZN(n58) );
  OR2_X2 U335 ( .A1(B[10]), .A2(A[10]), .ZN(n411) );
  NAND3_X1 U525 ( .A1(n169), .A2(n170), .A3(n171), .ZN(n168) );
  NAND3_X1 U531 ( .A1(n197), .A2(net537591), .A3(n198), .ZN(n196) );
  NAND3_X1 U567 ( .A1(n60), .A2(n376), .A3(n506), .ZN(n398) );
  NAND3_X1 U574 ( .A1(n5), .A2(n80), .A3(n46), .ZN(n433) );
  NAND3_X1 U578 ( .A1(n418), .A2(n64), .A3(n1), .ZN(n443) );
  NAND3_X1 U579 ( .A1(n5), .A2(n80), .A3(n46), .ZN(n418) );
  NAND3_X1 U583 ( .A1(n320), .A2(n318), .A3(n279), .ZN(n72) );
  NAND3_X1 U585 ( .A1(A[2]), .A2(B[2]), .A3(n279), .ZN(n386) );
  OR2_X2 U18 ( .A1(B[21]), .A2(A[21]), .ZN(n326) );
  OR2_X2 U95 ( .A1(B[26]), .A2(A[26]), .ZN(net507345) );
  OAI21_X2 U231 ( .B1(n456), .B2(n538), .A(n269), .ZN(n284) );
  AND2_X1 U2 ( .A1(n290), .A2(n270), .ZN(n456) );
  OR2_X1 U3 ( .A1(B[8]), .A2(A[8]), .ZN(n57) );
  NOR2_X1 U5 ( .A1(B[13]), .A2(A[13]), .ZN(n44) );
  AND2_X1 U6 ( .A1(n448), .A2(n447), .ZN(SUM[0]) );
  INV_X1 U7 ( .A(n456), .ZN(n288) );
  OR2_X1 U8 ( .A1(B[17]), .A2(A[17]), .ZN(n350) );
  OR2_X1 U9 ( .A1(B[16]), .A2(A[16]), .ZN(n349) );
  OR2_X1 U10 ( .A1(B[18]), .A2(A[18]), .ZN(n341) );
  OR2_X1 U11 ( .A1(B[20]), .A2(A[20]), .ZN(net507383) );
  OR2_X1 U12 ( .A1(B[25]), .A2(A[25]), .ZN(net507343) );
  OR2_X1 U13 ( .A1(B[28]), .A2(A[28]), .ZN(net507306) );
  OR2_X1 U14 ( .A1(B[29]), .A2(A[29]), .ZN(net507307) );
  OR2_X1 U15 ( .A1(B[40]), .A2(A[40]), .ZN(n248) );
  OR2_X1 U16 ( .A1(B[41]), .A2(A[41]), .ZN(n242) );
  OR2_X1 U17 ( .A1(B[42]), .A2(A[42]), .ZN(n243) );
  OR2_X1 U19 ( .A1(B[30]), .A2(A[30]), .ZN(net507290) );
  OR2_X1 U20 ( .A1(B[32]), .A2(A[32]), .ZN(n292) );
  OR2_X1 U21 ( .A1(B[33]), .A2(A[33]), .ZN(n293) );
  OR2_X1 U22 ( .A1(B[34]), .A2(A[34]), .ZN(n294) );
  OR2_X1 U23 ( .A1(B[45]), .A2(A[45]), .ZN(n223) );
  OR2_X1 U24 ( .A1(B[44]), .A2(A[44]), .ZN(n222) );
  OR2_X1 U25 ( .A1(B[46]), .A2(A[46]), .ZN(n209) );
  OR2_X1 U26 ( .A1(B[50]), .A2(A[50]), .ZN(n174) );
  OR2_X1 U27 ( .A1(B[48]), .A2(A[48]), .ZN(n172) );
  OR2_X1 U28 ( .A1(B[49]), .A2(A[49]), .ZN(n173) );
  OR2_X1 U29 ( .A1(B[52]), .A2(A[52]), .ZN(n153) );
  OR2_X1 U30 ( .A1(B[54]), .A2(A[54]), .ZN(n152) );
  OR2_X1 U31 ( .A1(B[53]), .A2(A[53]), .ZN(n154) );
  CLKBUF_X1 U32 ( .A(A[5]), .Z(n451) );
  AND2_X1 U33 ( .A1(n267), .A2(n271), .ZN(n452) );
  CLKBUF_X1 U34 ( .A(net507348), .Z(n453) );
  CLKBUF_X1 U35 ( .A(n247), .Z(n454) );
  INV_X1 U36 ( .A(n459), .ZN(n376) );
  NOR2_X1 U37 ( .A1(A[12]), .A2(B[12]), .ZN(n459) );
  INV_X1 U38 ( .A(n500), .ZN(n455) );
  AOI21_X1 U39 ( .B1(n351), .B2(n10), .A(net507300), .ZN(net538645) );
  OR2_X1 U40 ( .A1(B[14]), .A2(A[14]), .ZN(n369) );
  AND2_X1 U41 ( .A1(net507336), .A2(net507295), .ZN(net537128) );
  OR2_X2 U42 ( .A1(A[23]), .A2(B[23]), .ZN(n323) );
  INV_X1 U43 ( .A(n558), .ZN(n457) );
  OAI21_X1 U44 ( .B1(n339), .B2(n338), .A(n340), .ZN(net507300) );
  OAI21_X1 U45 ( .B1(n13), .B2(n322), .A(n323), .ZN(n458) );
  OAI21_X1 U46 ( .B1(n13), .B2(n322), .A(n323), .ZN(net507296) );
  CLKBUF_X1 U47 ( .A(n434), .Z(n460) );
  BUF_X1 U48 ( .A(n328), .Z(n461) );
  OR2_X1 U49 ( .A1(A[22]), .A2(B[22]), .ZN(n328) );
  OR2_X1 U50 ( .A1(n314), .A2(n515), .ZN(n462) );
  NAND2_X1 U51 ( .A1(n462), .A2(net535421), .ZN(net507279) );
  XNOR2_X1 U52 ( .A(n19), .B(n463), .ZN(SUM[8]) );
  NAND2_X1 U53 ( .A1(n57), .A2(n62), .ZN(n463) );
  INV_X1 U54 ( .A(n466), .ZN(n201) );
  OR2_X1 U55 ( .A1(B[43]), .A2(A[43]), .ZN(n238) );
  AND4_X1 U56 ( .A1(net507306), .A2(net507307), .A3(net507290), .A4(net507291), 
        .ZN(net535421) );
  OAI21_X1 U57 ( .B1(n555), .B2(n504), .A(n467), .ZN(n464) );
  CLKBUF_X1 U58 ( .A(n202), .Z(n465) );
  AND4_X1 U59 ( .A1(n248), .A2(n242), .A3(n243), .A4(n238), .ZN(n466) );
  CLKBUF_X1 U60 ( .A(n407), .Z(n467) );
  NAND3_X1 U61 ( .A1(n263), .A2(n268), .A3(n452), .ZN(n202) );
  OR2_X1 U62 ( .A1(B[36]), .A2(A[36]), .ZN(n271) );
  OR2_X1 U63 ( .A1(B[37]), .A2(A[37]), .ZN(n267) );
  OR2_X1 U64 ( .A1(B[38]), .A2(A[38]), .ZN(n268) );
  AND2_X1 U65 ( .A1(n312), .A2(n301), .ZN(n468) );
  OAI21_X1 U66 ( .B1(net537128), .B2(n512), .A(net507285), .ZN(n469) );
  XNOR2_X1 U67 ( .A(n470), .B(n471), .ZN(SUM[9]) );
  NOR2_X1 U68 ( .A1(n52), .A2(n53), .ZN(n470) );
  NOR2_X1 U69 ( .A1(n8), .A2(n505), .ZN(n471) );
  OR2_X1 U70 ( .A1(B[9]), .A2(A[9]), .ZN(n419) );
  OAI21_X1 U72 ( .B1(n542), .B2(n488), .A(n244), .ZN(n472) );
  OAI21_X1 U73 ( .B1(n488), .B2(n542), .A(n244), .ZN(n252) );
  XNOR2_X1 U74 ( .A(n473), .B(net537591), .ZN(SUM[32]) );
  NAND2_X1 U75 ( .A1(n292), .A2(n301), .ZN(n473) );
  XOR2_X1 U76 ( .A(n33), .B(n474), .Z(SUM[34]) );
  AND2_X1 U77 ( .A1(n294), .A2(n303), .ZN(n474) );
  XOR2_X1 U78 ( .A(n475), .B(n158), .Z(SUM[54]) );
  AND2_X1 U79 ( .A1(n152), .A2(n149), .ZN(n475) );
  XOR2_X1 U80 ( .A(n476), .B(n162), .Z(SUM[53]) );
  AND2_X1 U81 ( .A1(n154), .A2(n148), .ZN(n476) );
  XOR2_X1 U82 ( .A(n486), .B(n477), .Z(SUM[25]) );
  NAND2_X1 U83 ( .A1(net507367), .A2(net507347), .ZN(n477) );
  XOR2_X1 U84 ( .A(net537128), .B(n478), .Z(SUM[28]) );
  NAND2_X1 U85 ( .A1(net507306), .A2(net507285), .ZN(n478) );
  XNOR2_X1 U86 ( .A(n479), .B(n480), .ZN(SUM[7]) );
  AND2_X1 U87 ( .A1(n63), .A2(n64), .ZN(n479) );
  AND2_X1 U88 ( .A1(n58), .A2(n434), .ZN(n480) );
  XOR2_X1 U89 ( .A(n500), .B(n481), .Z(SUM[20]) );
  AND2_X1 U90 ( .A1(net507383), .A2(net507382), .ZN(n481) );
  INV_X1 U91 ( .A(n387), .ZN(n563) );
  INV_X1 U92 ( .A(n20), .ZN(n489) );
  NOR2_X1 U93 ( .A1(net537590), .A2(n514), .ZN(n314) );
  INV_X1 U94 ( .A(net507295), .ZN(n515) );
  AOI21_X1 U96 ( .B1(n401), .B2(n400), .A(n551), .ZN(n31) );
  NOR2_X1 U97 ( .A1(n507), .A2(n505), .ZN(n439) );
  AND2_X1 U98 ( .A1(net507302), .A2(n10), .ZN(n16) );
  NOR2_X1 U99 ( .A1(n499), .A2(net507301), .ZN(net507302) );
  INV_X1 U100 ( .A(net537591), .ZN(n490) );
  NAND2_X1 U101 ( .A1(n382), .A2(n55), .ZN(n19) );
  NOR2_X1 U102 ( .A1(n507), .A2(n428), .ZN(n425) );
  INV_X1 U103 ( .A(n139), .ZN(n496) );
  INV_X1 U104 ( .A(n165), .ZN(n498) );
  INV_X1 U105 ( .A(n108), .ZN(n495) );
  INV_X1 U106 ( .A(n221), .ZN(n537) );
  OR2_X1 U107 ( .A1(net507301), .A2(n510), .ZN(net507297) );
  INV_X1 U108 ( .A(n129), .ZN(n561) );
  NAND2_X1 U109 ( .A1(n564), .A2(n73), .ZN(n387) );
  INV_X1 U110 ( .A(n72), .ZN(n564) );
  NOR2_X1 U111 ( .A1(n83), .A2(n527), .ZN(SUM[64]) );
  NAND2_X1 U112 ( .A1(n326), .A2(n329), .ZN(n336) );
  NAND2_X1 U113 ( .A1(n549), .A2(n374), .ZN(n396) );
  XOR2_X1 U115 ( .A(n482), .B(n454), .Z(SUM[40]) );
  AND2_X1 U116 ( .A1(n248), .A2(n245), .ZN(n482) );
  NAND2_X1 U117 ( .A1(n172), .A2(n180), .ZN(n194) );
  NAND2_X1 U118 ( .A1(n293), .A2(n302), .ZN(n311) );
  XOR2_X1 U119 ( .A(n483), .B(n469), .Z(SUM[29]) );
  AND2_X1 U120 ( .A1(net507307), .A2(net507286), .ZN(n483) );
  NAND2_X1 U121 ( .A1(n173), .A2(n182), .ZN(n192) );
  NAND2_X1 U122 ( .A1(n222), .A2(n213), .ZN(n234) );
  NAND2_X1 U123 ( .A1(n223), .A2(n214), .ZN(n231) );
  NAND2_X1 U124 ( .A1(n242), .A2(n244), .ZN(n257) );
  NAND2_X1 U125 ( .A1(n243), .A2(n240), .ZN(n253) );
  NAND2_X1 U126 ( .A1(n349), .A2(n348), .ZN(n361) );
  NAND2_X1 U127 ( .A1(net507340), .A2(net507341), .ZN(net507338) );
  NAND2_X1 U128 ( .A1(net507346), .A2(net507347), .ZN(net507344) );
  NAND2_X1 U130 ( .A1(n264), .A2(n265), .ZN(n262) );
  NOR2_X1 U131 ( .A1(n14), .A2(n266), .ZN(n261) );
  AND2_X1 U132 ( .A1(n269), .A2(n270), .ZN(n14) );
  NAND2_X1 U133 ( .A1(net507345), .A2(net507341), .ZN(net507360) );
  XOR2_X1 U134 ( .A(n356), .B(n484), .Z(SUM[18]) );
  AND2_X1 U135 ( .A1(n341), .A2(n345), .ZN(n484) );
  NOR2_X1 U136 ( .A1(n518), .A2(n517), .ZN(n321) );
  INV_X1 U137 ( .A(net507340), .ZN(n518) );
  INV_X1 U138 ( .A(net507383), .ZN(n546) );
  AND2_X1 U139 ( .A1(n326), .A2(net507383), .ZN(n17) );
  OAI21_X1 U140 ( .B1(n497), .B2(n525), .A(n148), .ZN(n158) );
  INV_X1 U141 ( .A(n162), .ZN(n497) );
  OAI21_X1 U142 ( .B1(n492), .B2(n533), .A(n117), .ZN(n132) );
  INV_X1 U143 ( .A(n136), .ZN(n492) );
  OAI21_X1 U144 ( .B1(n491), .B2(n521), .A(n182), .ZN(n186) );
  OAI21_X1 U145 ( .B1(n535), .B2(n498), .A(n147), .ZN(n162) );
  INV_X1 U146 ( .A(n153), .ZN(n535) );
  OAI21_X1 U147 ( .B1(n141), .B2(n498), .A(n143), .ZN(n139) );
  NAND4_X1 U148 ( .A1(n153), .A2(n154), .A3(n152), .A4(n155), .ZN(n141) );
  AOI21_X1 U149 ( .B1(n144), .B2(n145), .A(n47), .ZN(n143) );
  OAI211_X1 U150 ( .C1(n525), .C2(n147), .A(n148), .B(n149), .ZN(n145) );
  OAI21_X1 U151 ( .B1(n495), .B2(n529), .A(n94), .ZN(n105) );
  OAI21_X1 U152 ( .B1(n494), .B2(n528), .A(n93), .ZN(n101) );
  INV_X1 U153 ( .A(n105), .ZN(n494) );
  OAI21_X1 U154 ( .B1(n534), .B2(n496), .A(n116), .ZN(n136) );
  INV_X1 U155 ( .A(n122), .ZN(n534) );
  OAI21_X1 U156 ( .B1(n110), .B2(n496), .A(n112), .ZN(n108) );
  NAND4_X1 U157 ( .A1(n122), .A2(n123), .A3(n121), .A4(n124), .ZN(n110) );
  AOI21_X1 U158 ( .B1(n113), .B2(n114), .A(n48), .ZN(n112) );
  OAI211_X1 U159 ( .C1(n533), .C2(n116), .A(n117), .B(n118), .ZN(n114) );
  NAND2_X1 U160 ( .A1(net507290), .A2(net507287), .ZN(net507318) );
  NAND2_X1 U161 ( .A1(n461), .A2(n325), .ZN(n334) );
  OAI21_X1 U162 ( .B1(n358), .B2(n511), .A(n346), .ZN(n356) );
  NAND2_X1 U163 ( .A1(n29), .A2(net507291), .ZN(net507312) );
  OAI21_X1 U164 ( .B1(n487), .B2(n541), .A(n214), .ZN(n227) );
  XNOR2_X1 U165 ( .A(n20), .B(n291), .ZN(SUM[36]) );
  NAND2_X1 U166 ( .A1(n271), .A2(n270), .ZN(n291) );
  NOR2_X1 U167 ( .A1(n509), .A2(n511), .ZN(n359) );
  INV_X1 U168 ( .A(n346), .ZN(n509) );
  NOR2_X1 U169 ( .A1(n555), .A2(n11), .ZN(n423) );
  XNOR2_X1 U170 ( .A(n453), .B(net507370), .ZN(SUM[24]) );
  NAND2_X1 U171 ( .A1(net507349), .A2(net507347), .ZN(net507370) );
  XOR2_X1 U172 ( .A(n485), .B(n288), .Z(SUM[37]) );
  AND2_X1 U173 ( .A1(n267), .A2(n269), .ZN(n485) );
  XNOR2_X1 U174 ( .A(n166), .B(n165), .ZN(SUM[52]) );
  NAND2_X1 U175 ( .A1(n153), .A2(n147), .ZN(n166) );
  XNOR2_X1 U176 ( .A(n285), .B(n284), .ZN(SUM[38]) );
  NAND2_X1 U177 ( .A1(n268), .A2(n265), .ZN(n285) );
  XNOR2_X1 U178 ( .A(n187), .B(n186), .ZN(SUM[50]) );
  NAND2_X1 U179 ( .A1(n174), .A2(n181), .ZN(n187) );
  XNOR2_X1 U180 ( .A(n228), .B(n227), .ZN(SUM[46]) );
  NAND2_X1 U181 ( .A1(n209), .A2(n215), .ZN(n228) );
  XNOR2_X1 U182 ( .A(n140), .B(n139), .ZN(SUM[56]) );
  NAND2_X1 U183 ( .A1(n122), .A2(n116), .ZN(n140) );
  XNOR2_X1 U184 ( .A(n137), .B(n136), .ZN(SUM[57]) );
  NAND2_X1 U185 ( .A1(n123), .A2(n117), .ZN(n137) );
  XNOR2_X1 U186 ( .A(n134), .B(n132), .ZN(SUM[58]) );
  NAND2_X1 U187 ( .A1(n121), .A2(n118), .ZN(n134) );
  XNOR2_X1 U188 ( .A(n109), .B(n108), .ZN(SUM[60]) );
  NAND2_X1 U189 ( .A1(n107), .A2(n94), .ZN(n109) );
  XNOR2_X1 U190 ( .A(n106), .B(n105), .ZN(SUM[61]) );
  NAND2_X1 U191 ( .A1(n104), .A2(n93), .ZN(n106) );
  XNOR2_X1 U192 ( .A(n102), .B(n101), .ZN(SUM[62]) );
  NAND2_X1 U193 ( .A1(n100), .A2(n90), .ZN(n102) );
  OAI21_X1 U194 ( .B1(n544), .B2(n468), .A(n302), .ZN(n33) );
  XNOR2_X1 U195 ( .A(n97), .B(n98), .ZN(SUM[63]) );
  NAND2_X1 U196 ( .A1(n89), .A2(n85), .ZN(n97) );
  OAI21_X1 U197 ( .B1(n493), .B2(n526), .A(n90), .ZN(n98) );
  INV_X1 U198 ( .A(n101), .ZN(n493) );
  XNOR2_X1 U199 ( .A(n331), .B(n330), .ZN(SUM[23]) );
  NAND2_X1 U200 ( .A1(n324), .A2(n323), .ZN(n330) );
  NAND2_X1 U201 ( .A1(n332), .A2(n325), .ZN(n331) );
  XNOR2_X1 U202 ( .A(n436), .B(n437), .ZN(SUM[10]) );
  NOR2_X1 U203 ( .A1(n552), .A2(n553), .ZN(n437) );
  AOI21_X1 U204 ( .B1(n440), .B2(n439), .A(n8), .ZN(n436) );
  INV_X1 U205 ( .A(n411), .ZN(n553) );
  INV_X1 U206 ( .A(n374), .ZN(n550) );
  OAI21_X1 U207 ( .B1(n236), .B2(n237), .A(n238), .ZN(n217) );
  NAND2_X1 U208 ( .A1(n239), .A2(n240), .ZN(n237) );
  NOR2_X1 U209 ( .A1(n15), .A2(n241), .ZN(n236) );
  AND2_X1 U210 ( .A1(n244), .A2(n245), .ZN(n15) );
  NOR2_X1 U211 ( .A1(n343), .A2(n344), .ZN(n338) );
  NAND2_X1 U212 ( .A1(n345), .A2(n346), .ZN(n344) );
  OAI21_X1 U213 ( .B1(net537128), .B2(n512), .A(net507285), .ZN(n26) );
  INV_X1 U214 ( .A(net507306), .ZN(n512) );
  NAND2_X1 U215 ( .A1(net507282), .A2(net507283), .ZN(net507280) );
  AND2_X1 U216 ( .A1(net507291), .A2(net507290), .ZN(net507282) );
  OAI211_X1 U217 ( .C1(n513), .C2(net507285), .A(net507286), .B(net507287), 
        .ZN(net507283) );
  NOR2_X1 U218 ( .A1(n561), .A2(n69), .ZN(n77) );
  XNOR2_X1 U219 ( .A(n388), .B(n389), .ZN(SUM[15]) );
  NAND2_X1 U220 ( .A1(n368), .A2(n9), .ZN(n389) );
  OAI21_X1 U221 ( .B1(n390), .B2(n391), .A(n373), .ZN(n388) );
  NAND2_X1 U222 ( .A1(n549), .A2(n369), .ZN(n391) );
  XNOR2_X1 U223 ( .A(n156), .B(n157), .ZN(SUM[55]) );
  NOR2_X1 U224 ( .A1(n522), .A2(n47), .ZN(n157) );
  AOI21_X1 U225 ( .B1(n152), .B2(n158), .A(n524), .ZN(n156) );
  INV_X1 U226 ( .A(n149), .ZN(n524) );
  XNOR2_X1 U227 ( .A(n130), .B(n131), .ZN(SUM[59]) );
  NOR2_X1 U228 ( .A1(n530), .A2(n48), .ZN(n131) );
  AOI21_X1 U229 ( .B1(n121), .B2(n132), .A(n532), .ZN(n130) );
  INV_X1 U230 ( .A(n118), .ZN(n532) );
  AND2_X1 U232 ( .A1(net507343), .A2(net507346), .ZN(n486) );
  XNOR2_X1 U233 ( .A(n250), .B(n249), .ZN(SUM[43]) );
  NAND2_X1 U234 ( .A1(n239), .A2(n238), .ZN(n249) );
  XNOR2_X1 U235 ( .A(n183), .B(n184), .ZN(SUM[51]) );
  NAND2_X1 U236 ( .A1(n175), .A2(n178), .ZN(n183) );
  NAND2_X1 U237 ( .A1(n181), .A2(n185), .ZN(n184) );
  NAND2_X1 U238 ( .A1(n174), .A2(n186), .ZN(n185) );
  OAI21_X1 U239 ( .B1(n504), .B2(n555), .A(n467), .ZN(n380) );
  NAND2_X1 U240 ( .A1(n417), .A2(n64), .ZN(n431) );
  NAND4_X1 U241 ( .A1(n369), .A2(n549), .A3(n376), .A4(n9), .ZN(n363) );
  AOI21_X1 U242 ( .B1(n508), .B2(n55), .A(n56), .ZN(n53) );
  XNOR2_X1 U243 ( .A(n404), .B(n405), .ZN(SUM[12]) );
  NAND2_X1 U244 ( .A1(n376), .A2(n375), .ZN(n404) );
  NAND2_X1 U245 ( .A1(n506), .A2(n19), .ZN(n406) );
  NOR2_X1 U246 ( .A1(n503), .A2(n378), .ZN(n362) );
  OAI21_X1 U247 ( .B1(n563), .B2(n385), .A(n18), .ZN(n381) );
  NOR2_X1 U248 ( .A1(n44), .A2(n375), .ZN(n371) );
  OAI21_X1 U249 ( .B1(n216), .B2(n201), .A(n217), .ZN(n204) );
  AOI21_X1 U250 ( .B1(n536), .B2(n219), .A(n537), .ZN(n216) );
  OAI21_X1 U251 ( .B1(n543), .B2(n297), .A(n298), .ZN(n219) );
  NOR2_X1 U252 ( .A1(n511), .A2(n348), .ZN(n343) );
  NOR2_X1 U253 ( .A1(n522), .A2(n523), .ZN(n144) );
  INV_X1 U254 ( .A(n152), .ZN(n523) );
  NOR2_X1 U255 ( .A1(n530), .A2(n531), .ZN(n113) );
  INV_X1 U256 ( .A(n121), .ZN(n531) );
  NAND2_X1 U257 ( .A1(n167), .A2(n168), .ZN(n165) );
  AOI21_X1 U258 ( .B1(n169), .B2(n176), .A(n520), .ZN(n167) );
  OAI211_X1 U259 ( .C1(n521), .C2(n180), .A(n181), .B(n182), .ZN(n176) );
  INV_X1 U260 ( .A(n350), .ZN(n511) );
  OAI21_X1 U261 ( .B1(n428), .B2(n414), .A(n429), .ZN(n427) );
  OAI21_X1 U262 ( .B1(n366), .B2(n367), .A(n368), .ZN(n365) );
  NAND2_X1 U263 ( .A1(n369), .A2(n370), .ZN(n367) );
  NOR2_X1 U264 ( .A1(n372), .A2(n371), .ZN(n366) );
  OAI21_X1 U265 ( .B1(n2), .B2(n516), .A(net507346), .ZN(net507358) );
  INV_X1 U266 ( .A(n44), .ZN(n549) );
  OAI21_X1 U267 ( .B1(n539), .B2(n207), .A(n208), .ZN(n205) );
  INV_X1 U268 ( .A(n211), .ZN(n539) );
  OAI211_X1 U269 ( .C1(n541), .C2(n213), .A(n214), .B(n215), .ZN(n211) );
  NAND2_X1 U270 ( .A1(n411), .A2(n419), .ZN(n428) );
  INV_X1 U271 ( .A(n293), .ZN(n544) );
  XNOR2_X1 U272 ( .A(n395), .B(n394), .ZN(SUM[14]) );
  NAND2_X1 U273 ( .A1(n373), .A2(n369), .ZN(n394) );
  OAI21_X1 U274 ( .B1(n39), .B2(n44), .A(n374), .ZN(n395) );
  INV_X1 U275 ( .A(n299), .ZN(n543) );
  OAI211_X1 U276 ( .C1(n544), .C2(n301), .A(n302), .B(n303), .ZN(n299) );
  NAND2_X1 U277 ( .A1(n560), .A2(n554), .ZN(n407) );
  INV_X1 U278 ( .A(n409), .ZN(n555) );
  NAND2_X1 U279 ( .A1(n312), .A2(n301), .ZN(n310) );
  NAND2_X1 U280 ( .A1(n258), .A2(n245), .ZN(n256) );
  NAND2_X1 U281 ( .A1(n193), .A2(n180), .ZN(n189) );
  INV_X1 U282 ( .A(n419), .ZN(n505) );
  INV_X1 U283 ( .A(n57), .ZN(n507) );
  INV_X1 U284 ( .A(net507307), .ZN(n513) );
  INV_X1 U285 ( .A(n104), .ZN(n528) );
  INV_X1 U286 ( .A(n100), .ZN(n526) );
  INV_X1 U287 ( .A(n155), .ZN(n522) );
  INV_X1 U288 ( .A(n124), .ZN(n530) );
  INV_X1 U289 ( .A(n267), .ZN(n538) );
  INV_X1 U290 ( .A(n107), .ZN(n529) );
  INV_X1 U291 ( .A(n154), .ZN(n525) );
  INV_X1 U292 ( .A(n123), .ZN(n533) );
  INV_X1 U293 ( .A(n173), .ZN(n521) );
  INV_X1 U294 ( .A(n223), .ZN(n541) );
  NAND2_X1 U295 ( .A1(n373), .A2(n374), .ZN(n372) );
  AND4_X1 U296 ( .A1(n6), .A2(n350), .A3(n341), .A4(n349), .ZN(n10) );
  AND2_X1 U297 ( .A1(n560), .A2(n554), .ZN(n11) );
  INV_X1 U298 ( .A(n375), .ZN(n551) );
  AND2_X1 U299 ( .A1(n174), .A2(n175), .ZN(n169) );
  INV_X1 U300 ( .A(n242), .ZN(n542) );
  NAND2_X1 U301 ( .A1(n242), .A2(n243), .ZN(n241) );
  NAND2_X1 U302 ( .A1(n324), .A2(n325), .ZN(n322) );
  AND3_X1 U303 ( .A1(n326), .A2(n327), .A3(n328), .ZN(n13) );
  NAND2_X1 U304 ( .A1(n329), .A2(net507382), .ZN(n327) );
  NAND2_X1 U305 ( .A1(n267), .A2(n268), .ZN(n266) );
  INV_X1 U306 ( .A(net507343), .ZN(n516) );
  INV_X1 U307 ( .A(n429), .ZN(n552) );
  INV_X1 U308 ( .A(n348), .ZN(n545) );
  NAND2_X1 U309 ( .A1(n6), .A2(n340), .ZN(n353) );
  NAND2_X1 U310 ( .A1(n356), .A2(n341), .ZN(n355) );
  INV_X1 U311 ( .A(n326), .ZN(n547) );
  INV_X1 U312 ( .A(n64), .ZN(n557) );
  INV_X1 U313 ( .A(n178), .ZN(n520) );
  INV_X1 U314 ( .A(net507341), .ZN(n519) );
  AND2_X1 U315 ( .A1(n172), .A2(n173), .ZN(n170) );
  XNOR2_X1 U316 ( .A(n125), .B(n126), .ZN(SUM[5]) );
  AOI21_X1 U317 ( .B1(n129), .B2(n82), .A(n46), .ZN(n125) );
  NOR2_X1 U318 ( .A1(n444), .A2(n558), .ZN(n126) );
  XNOR2_X1 U320 ( .A(n273), .B(n274), .ZN(SUM[3]) );
  OAI21_X1 U321 ( .B1(n566), .B2(n565), .A(n277), .ZN(n274) );
  NAND2_X1 U322 ( .A1(n279), .A2(n280), .ZN(n273) );
  INV_X1 U323 ( .A(n278), .ZN(n566) );
  XNOR2_X1 U324 ( .A(n352), .B(n568), .ZN(SUM[1]) );
  NAND2_X1 U325 ( .A1(n318), .A2(n317), .ZN(n352) );
  XNOR2_X1 U326 ( .A(n315), .B(n278), .ZN(SUM[2]) );
  NAND2_X1 U327 ( .A1(n320), .A2(n277), .ZN(n315) );
  XNOR2_X1 U328 ( .A(n561), .B(n190), .ZN(SUM[4]) );
  NOR2_X1 U329 ( .A1(n559), .A2(n46), .ZN(n190) );
  INV_X1 U330 ( .A(n80), .ZN(n558) );
  INV_X1 U331 ( .A(n82), .ZN(n559) );
  AOI21_X1 U332 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  NAND2_X1 U333 ( .A1(n89), .A2(n90), .ZN(n88) );
  NOR2_X1 U334 ( .A1(n526), .A2(n528), .ZN(n86) );
  OAI211_X1 U336 ( .C1(n495), .C2(n529), .A(n93), .B(n94), .ZN(n87) );
  NAND2_X1 U337 ( .A1(n562), .A2(n387), .ZN(n129) );
  INV_X1 U338 ( .A(n385), .ZN(n562) );
  NAND2_X1 U339 ( .A1(n129), .A2(n415), .ZN(n55) );
  NOR2_X1 U340 ( .A1(n558), .A2(n559), .ZN(n416) );
  NAND2_X1 U341 ( .A1(n316), .A2(n317), .ZN(n278) );
  NAND2_X1 U342 ( .A1(n318), .A2(n568), .ZN(n316) );
  NAND2_X1 U343 ( .A1(n82), .A2(n80), .ZN(n69) );
  NAND2_X1 U344 ( .A1(n447), .A2(n317), .ZN(n73) );
  INV_X1 U345 ( .A(n447), .ZN(n568) );
  NOR2_X1 U346 ( .A1(n68), .A2(n69), .ZN(n65) );
  NOR2_X1 U347 ( .A1(n385), .A2(n70), .ZN(n68) );
  NOR2_X1 U348 ( .A1(n567), .A2(n72), .ZN(n70) );
  INV_X1 U349 ( .A(n73), .ZN(n567) );
  INV_X1 U350 ( .A(n320), .ZN(n565) );
  INV_X1 U351 ( .A(n85), .ZN(n527) );
  OAI21_X1 U352 ( .B1(n413), .B2(n62), .A(n414), .ZN(n410) );
  NAND2_X1 U353 ( .A1(B[13]), .A2(A[13]), .ZN(n374) );
  NAND2_X1 U354 ( .A1(A[6]), .A2(B[6]), .ZN(n64) );
  NAND2_X1 U355 ( .A1(B[33]), .A2(A[33]), .ZN(n302) );
  NAND2_X1 U356 ( .A1(A[8]), .A2(B[8]), .ZN(n62) );
  OR2_X1 U357 ( .A1(B[58]), .A2(A[58]), .ZN(n121) );
  NAND2_X1 U358 ( .A1(A[22]), .A2(B[22]), .ZN(n325) );
  NAND2_X1 U359 ( .A1(A[12]), .A2(B[12]), .ZN(n375) );
  NAND2_X1 U360 ( .A1(B[29]), .A2(A[29]), .ZN(net507286) );
  NAND2_X1 U361 ( .A1(B[21]), .A2(A[21]), .ZN(n329) );
  NOR2_X1 U362 ( .A1(B[6]), .A2(A[6]), .ZN(n34) );
  NAND2_X1 U363 ( .A1(B[26]), .A2(A[26]), .ZN(net507341) );
  NAND2_X1 U364 ( .A1(B[32]), .A2(A[32]), .ZN(n301) );
  NAND2_X1 U365 ( .A1(B[24]), .A2(A[24]), .ZN(net507347) );
  NAND2_X1 U366 ( .A1(B[48]), .A2(A[48]), .ZN(n180) );
  NAND2_X1 U367 ( .A1(B[28]), .A2(A[28]), .ZN(net507285) );
  NAND2_X1 U368 ( .A1(B[62]), .A2(A[62]), .ZN(n90) );
  NAND2_X1 U369 ( .A1(B[16]), .A2(A[16]), .ZN(n348) );
  NAND2_X1 U370 ( .A1(B[61]), .A2(A[61]), .ZN(n93) );
  NAND2_X1 U371 ( .A1(B[53]), .A2(A[53]), .ZN(n148) );
  NAND2_X1 U372 ( .A1(B[57]), .A2(A[57]), .ZN(n117) );
  NAND2_X1 U373 ( .A1(B[45]), .A2(A[45]), .ZN(n214) );
  NAND2_X1 U374 ( .A1(B[54]), .A2(A[54]), .ZN(n149) );
  NAND2_X1 U375 ( .A1(B[58]), .A2(A[58]), .ZN(n118) );
  NAND2_X1 U376 ( .A1(B[17]), .A2(A[17]), .ZN(n346) );
  NAND2_X1 U377 ( .A1(B[52]), .A2(A[52]), .ZN(n147) );
  NAND2_X1 U378 ( .A1(B[56]), .A2(A[56]), .ZN(n116) );
  NAND2_X1 U379 ( .A1(B[49]), .A2(A[49]), .ZN(n182) );
  NAND2_X1 U380 ( .A1(B[60]), .A2(A[60]), .ZN(n94) );
  NAND2_X1 U381 ( .A1(B[50]), .A2(A[50]), .ZN(n181) );
  NAND2_X1 U382 ( .A1(A[14]), .A2(B[14]), .ZN(n373) );
  NAND2_X1 U383 ( .A1(B[38]), .A2(A[38]), .ZN(n265) );
  NAND2_X1 U384 ( .A1(B[37]), .A2(A[37]), .ZN(n269) );
  NAND2_X1 U385 ( .A1(B[34]), .A2(A[34]), .ZN(n303) );
  NAND2_X1 U386 ( .A1(B[40]), .A2(A[40]), .ZN(n245) );
  NAND2_X1 U387 ( .A1(B[20]), .A2(A[20]), .ZN(net507382) );
  NAND2_X1 U388 ( .A1(B[42]), .A2(A[42]), .ZN(n240) );
  NAND2_X1 U389 ( .A1(B[46]), .A2(A[46]), .ZN(n215) );
  NAND2_X1 U390 ( .A1(B[44]), .A2(A[44]), .ZN(n213) );
  NAND2_X1 U391 ( .A1(B[41]), .A2(A[41]), .ZN(n244) );
  NAND2_X1 U392 ( .A1(B[30]), .A2(A[30]), .ZN(net507287) );
  OR2_X1 U393 ( .A1(B[57]), .A2(A[57]), .ZN(n123) );
  NAND2_X1 U394 ( .A1(A[15]), .A2(B[15]), .ZN(n368) );
  OR2_X1 U395 ( .A1(B[56]), .A2(A[56]), .ZN(n122) );
  NAND2_X1 U396 ( .A1(A[10]), .A2(B[10]), .ZN(n429) );
  NAND2_X1 U397 ( .A1(B[36]), .A2(A[36]), .ZN(n270) );
  NAND2_X1 U398 ( .A1(B[51]), .A2(A[51]), .ZN(n178) );
  NAND2_X1 U399 ( .A1(B[63]), .A2(A[63]), .ZN(n89) );
  OR2_X1 U400 ( .A1(B[15]), .A2(A[15]), .ZN(n9) );
  AND2_X1 U401 ( .A1(B[55]), .A2(A[55]), .ZN(n47) );
  AND2_X1 U402 ( .A1(B[59]), .A2(A[59]), .ZN(n48) );
  OR2_X1 U403 ( .A1(A[31]), .A2(B[31]), .ZN(net507291) );
  OR2_X1 U404 ( .A1(B[55]), .A2(A[55]), .ZN(n155) );
  OR2_X1 U405 ( .A1(B[59]), .A2(A[59]), .ZN(n124) );
  OR2_X1 U406 ( .A1(B[24]), .A2(A[24]), .ZN(net507349) );
  OR2_X1 U407 ( .A1(B[63]), .A2(A[63]), .ZN(n85) );
  AND2_X1 U408 ( .A1(A[8]), .A2(B[8]), .ZN(n52) );
  OR2_X1 U409 ( .A1(B[60]), .A2(A[60]), .ZN(n107) );
  OR2_X1 U410 ( .A1(B[61]), .A2(A[61]), .ZN(n104) );
  OR2_X1 U411 ( .A1(B[62]), .A2(A[62]), .ZN(n100) );
  INV_X1 U412 ( .A(B[11]), .ZN(n560) );
  OR2_X1 U413 ( .A1(A[39]), .A2(B[39]), .ZN(n263) );
  OR2_X1 U414 ( .A1(B[47]), .A2(A[47]), .ZN(n210) );
  OR2_X1 U415 ( .A1(B[51]), .A2(A[51]), .ZN(n175) );
  AND2_X1 U416 ( .A1(n41), .A2(n80), .ZN(n66) );
  NAND2_X1 U417 ( .A1(B[4]), .A2(A[4]), .ZN(n78) );
  OR2_X1 U418 ( .A1(A[6]), .A2(B[6]), .ZN(n67) );
  OR2_X1 U419 ( .A1(A[6]), .A2(B[6]), .ZN(n5) );
  OR2_X1 U420 ( .A1(B[15]), .A2(A[15]), .ZN(n370) );
  OR2_X1 U421 ( .A1(B[4]), .A2(A[4]), .ZN(n82) );
  OR2_X1 U422 ( .A1(B[2]), .A2(A[2]), .ZN(n320) );
  OR2_X1 U423 ( .A1(B[1]), .A2(A[1]), .ZN(n318) );
  OR2_X1 U424 ( .A1(B[3]), .A2(A[3]), .ZN(n279) );
  OR2_X1 U425 ( .A1(B[0]), .A2(A[0]), .ZN(n448) );
  NAND2_X1 U426 ( .A1(B[1]), .A2(A[1]), .ZN(n317) );
  NAND2_X1 U427 ( .A1(n386), .A2(n280), .ZN(n385) );
  NAND2_X1 U428 ( .A1(B[0]), .A2(A[0]), .ZN(n447) );
  NAND2_X1 U429 ( .A1(B[2]), .A2(A[2]), .ZN(n277) );
  NAND2_X1 U430 ( .A1(B[3]), .A2(A[3]), .ZN(n280) );
  XNOR2_X1 U431 ( .A(n74), .B(n75), .ZN(SUM[6]) );
  NOR2_X1 U432 ( .A1(n77), .A2(n66), .ZN(n74) );
  XNOR2_X1 U433 ( .A(n392), .B(n396), .ZN(SUM[13]) );
  NOR2_X1 U434 ( .A1(n392), .A2(n550), .ZN(n390) );
  OAI21_X1 U435 ( .B1(n363), .B2(n362), .A(n548), .ZN(net537652) );
  NAND2_X1 U436 ( .A1(B[7]), .A2(A[7]), .ZN(n434) );
  NAND2_X1 U437 ( .A1(n58), .A2(n45), .ZN(n441) );
  OAI21_X1 U438 ( .B1(n431), .B2(n432), .A(n58), .ZN(n430) );
  AOI21_X1 U439 ( .B1(n58), .B2(n443), .A(n52), .ZN(n442) );
  NAND2_X1 U440 ( .A1(n57), .A2(n58), .ZN(n56) );
  AND3_X1 U441 ( .A1(n416), .A2(n556), .A3(n58), .ZN(n415) );
  AND3_X1 U442 ( .A1(n457), .A2(n82), .A3(n556), .ZN(n45) );
  AND4_X1 U443 ( .A1(n82), .A2(n80), .A3(n556), .A4(n58), .ZN(n18) );
  OAI21_X1 U444 ( .B1(n65), .B2(n66), .A(n556), .ZN(n63) );
  NAND2_X1 U445 ( .A1(n283), .A2(n265), .ZN(n282) );
  INV_X1 U446 ( .A(n380), .ZN(n503) );
  NAND2_X1 U447 ( .A1(n406), .A2(n464), .ZN(n405) );
  AND2_X1 U448 ( .A1(A[9]), .A2(B[9]), .ZN(n8) );
  AOI21_X1 U449 ( .B1(n410), .B2(n411), .A(n552), .ZN(n408) );
  NOR2_X1 U450 ( .A1(A[9]), .A2(B[9]), .ZN(n413) );
  NAND2_X1 U451 ( .A1(A[9]), .A2(B[9]), .ZN(n414) );
  NAND2_X1 U452 ( .A1(n268), .A2(n284), .ZN(n283) );
  AOI21_X1 U453 ( .B1(n540), .B2(n204), .A(n205), .ZN(n195) );
  NAND2_X1 U454 ( .A1(n333), .A2(n461), .ZN(n332) );
  NAND2_X1 U455 ( .A1(B[18]), .A2(A[18]), .ZN(n345) );
  AOI21_X1 U456 ( .B1(n401), .B2(n400), .A(n551), .ZN(n397) );
  OAI211_X1 U457 ( .C1(n561), .C2(n441), .A(n460), .B(n442), .ZN(n440) );
  NAND2_X1 U458 ( .A1(n433), .A2(n434), .ZN(n432) );
  NAND4_X1 U459 ( .A1(n1), .A2(n418), .A3(n434), .A4(n64), .ZN(n59) );
  NAND2_X1 U460 ( .A1(B[25]), .A2(A[25]), .ZN(net507346) );
  AND3_X1 U461 ( .A1(net507343), .A2(net507344), .A3(net507345), .ZN(n12) );
  NAND2_X1 U462 ( .A1(A[23]), .A2(B[23]), .ZN(n324) );
  XNOR2_X1 U463 ( .A(n192), .B(n189), .ZN(SUM[49]) );
  INV_X1 U464 ( .A(n189), .ZN(n491) );
  AND2_X1 U465 ( .A1(n398), .A2(n31), .ZN(n39) );
  NAND2_X1 U466 ( .A1(n398), .A2(n397), .ZN(n392) );
  NAND2_X1 U467 ( .A1(A[11]), .A2(B[11]), .ZN(n409) );
  INV_X1 U468 ( .A(A[11]), .ZN(n554) );
  XNOR2_X1 U469 ( .A(net507313), .B(net507312), .ZN(SUM[31]) );
  NAND2_X1 U470 ( .A1(net507287), .A2(net507314), .ZN(net507313) );
  NAND2_X1 U471 ( .A1(n251), .A2(n240), .ZN(n250) );
  AOI21_X1 U472 ( .B1(net507358), .B2(net507345), .A(n519), .ZN(net507352) );
  NAND2_X1 U473 ( .A1(B[31]), .A2(A[31]), .ZN(n29) );
  XNOR2_X1 U474 ( .A(n194), .B(n171), .ZN(SUM[48]) );
  NAND2_X1 U475 ( .A1(n171), .A2(n172), .ZN(n193) );
  NAND2_X1 U476 ( .A1(n195), .A2(n196), .ZN(n171) );
  XNOR2_X1 U477 ( .A(n334), .B(n40), .ZN(SUM[22]) );
  NAND2_X1 U478 ( .A1(n342), .A2(n341), .ZN(n339) );
  NAND2_X1 U479 ( .A1(B[43]), .A2(A[43]), .ZN(n239) );
  INV_X1 U480 ( .A(net537017), .ZN(n514) );
  NAND2_X1 U481 ( .A1(net507348), .A2(net537017), .ZN(net507336) );
  OR2_X1 U482 ( .A1(B[27]), .A2(A[27]), .ZN(net507339) );
  NOR2_X1 U483 ( .A1(n557), .A2(n34), .ZN(n75) );
  INV_X1 U484 ( .A(n34), .ZN(n556) );
  XNOR2_X1 U485 ( .A(n311), .B(n310), .ZN(SUM[33]) );
  NAND2_X1 U486 ( .A1(n382), .A2(n55), .ZN(n60) );
  XNOR2_X1 U487 ( .A(n354), .B(n353), .ZN(SUM[19]) );
  NAND2_X1 U488 ( .A1(n355), .A2(n345), .ZN(n354) );
  OAI21_X1 U489 ( .B1(n362), .B2(n363), .A(n548), .ZN(n351) );
  INV_X1 U490 ( .A(n365), .ZN(n548) );
  AOI21_X1 U491 ( .B1(n351), .B2(n349), .A(n545), .ZN(n358) );
  AOI21_X1 U492 ( .B1(n426), .B2(n425), .A(n427), .ZN(n422) );
  OAI211_X1 U493 ( .C1(n561), .C2(n441), .A(n62), .B(n430), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n422), .B(n423), .ZN(SUM[11]) );
  XNOR2_X1 U495 ( .A(n282), .B(n281), .ZN(SUM[39]) );
  INV_X1 U496 ( .A(net507339), .ZN(n517) );
  OAI21_X1 U497 ( .B1(n12), .B2(net507338), .A(net507339), .ZN(net507295) );
  AND4_X2 U498 ( .A1(net507349), .A2(net507343), .A3(net507345), .A4(net507339), .ZN(net537017) );
  NAND2_X1 U499 ( .A1(n208), .A2(n210), .ZN(n224) );
  NAND2_X1 U500 ( .A1(n209), .A2(n210), .ZN(n207) );
  NAND4_X1 U501 ( .A1(n222), .A2(n223), .A3(n209), .A4(n210), .ZN(n199) );
  XNOR2_X1 U502 ( .A(n257), .B(n256), .ZN(SUM[41]) );
  INV_X1 U503 ( .A(n256), .ZN(n488) );
  NAND2_X1 U504 ( .A1(n264), .A2(n263), .ZN(n281) );
  OAI21_X1 U505 ( .B1(n261), .B2(n262), .A(n263), .ZN(n221) );
  NOR2_X1 U506 ( .A1(n459), .A2(n11), .ZN(n400) );
  OAI21_X1 U507 ( .B1(n2), .B2(n516), .A(net507346), .ZN(n3) );
  AND2_X1 U508 ( .A1(net507367), .A2(net507347), .ZN(n2) );
  XNOR2_X1 U509 ( .A(net507360), .B(n3), .ZN(SUM[26]) );
  NAND2_X1 U510 ( .A1(net507122), .A2(n292), .ZN(n312) );
  XNOR2_X1 U511 ( .A(net507318), .B(net537206), .ZN(SUM[30]) );
  NAND2_X1 U512 ( .A1(A[27]), .A2(B[27]), .ZN(net507340) );
  OAI21_X1 U513 ( .B1(n547), .B2(n502), .A(n329), .ZN(n40) );
  OAI21_X1 U514 ( .B1(n502), .B2(n547), .A(n329), .ZN(n333) );
  INV_X1 U515 ( .A(n199), .ZN(n540) );
  NAND2_X1 U516 ( .A1(B[47]), .A2(A[47]), .ZN(n208) );
  XNOR2_X1 U517 ( .A(n231), .B(n230), .ZN(SUM[45]) );
  INV_X1 U518 ( .A(n230), .ZN(n487) );
  NAND2_X1 U519 ( .A1(n78), .A2(n79), .ZN(n41) );
  OAI21_X1 U520 ( .B1(n513), .B2(n501), .A(net507286), .ZN(net537206) );
  OAI21_X1 U521 ( .B1(n501), .B2(n513), .A(net507286), .ZN(n27) );
  NAND2_X1 U522 ( .A1(n59), .A2(n58), .ZN(n382) );
  INV_X1 U523 ( .A(n59), .ZN(n508) );
  NAND2_X1 U524 ( .A1(n232), .A2(n213), .ZN(n230) );
  NAND2_X1 U526 ( .A1(B[35]), .A2(A[35]), .ZN(n298) );
  OR2_X1 U527 ( .A1(B[35]), .A2(A[35]), .ZN(n295) );
  NAND2_X1 U528 ( .A1(n235), .A2(n217), .ZN(n233) );
  NAND2_X1 U529 ( .A1(n67), .A2(n444), .ZN(n417) );
  NAND2_X1 U530 ( .A1(n67), .A2(n444), .ZN(n1) );
  INV_X1 U532 ( .A(net507300), .ZN(n510) );
  XNOR2_X1 U533 ( .A(n36), .B(n359), .ZN(SUM[17]) );
  NAND2_X1 U534 ( .A1(net507290), .A2(n27), .ZN(net507314) );
  XNOR2_X1 U535 ( .A(net507352), .B(n321), .ZN(SUM[27]) );
  AND2_X1 U536 ( .A1(net507296), .A2(net507297), .ZN(net537590) );
  NAND2_X1 U537 ( .A1(n4), .A2(net507349), .ZN(net507367) );
  NAND2_X1 U538 ( .A1(A[39]), .A2(B[39]), .ZN(n264) );
  XNOR2_X1 U539 ( .A(n224), .B(n225), .ZN(SUM[47]) );
  NAND2_X1 U540 ( .A1(n226), .A2(n215), .ZN(n225) );
  INV_X1 U541 ( .A(net537652), .ZN(n499) );
  XNOR2_X1 U542 ( .A(net537652), .B(n361), .ZN(SUM[16]) );
  AOI21_X1 U543 ( .B1(net537652), .B2(n349), .A(n545), .ZN(n36) );
  NAND2_X1 U544 ( .A1(n408), .A2(n409), .ZN(n401) );
  INV_X1 U545 ( .A(n408), .ZN(n504) );
  OAI21_X1 U546 ( .B1(n455), .B2(net507301), .A(net507296), .ZN(net507348) );
  XNOR2_X1 U547 ( .A(net507395), .B(n336), .ZN(SUM[21]) );
  INV_X1 U548 ( .A(net538645), .ZN(n500) );
  OAI21_X1 U549 ( .B1(n455), .B2(net507301), .A(n458), .ZN(n4) );
  INV_X1 U550 ( .A(net507395), .ZN(n502) );
  OAI21_X1 U551 ( .B1(net538645), .B2(n546), .A(net507382), .ZN(net507395) );
  NAND2_X1 U552 ( .A1(A[19]), .A2(B[19]), .ZN(n340) );
  OR2_X1 U553 ( .A1(B[19]), .A2(A[19]), .ZN(n6) );
  OR2_X1 U554 ( .A1(A[19]), .A2(B[19]), .ZN(n342) );
  XNOR2_X1 U555 ( .A(n234), .B(n233), .ZN(SUM[44]) );
  NAND2_X1 U556 ( .A1(n233), .A2(n222), .ZN(n232) );
  AND2_X1 U557 ( .A1(n451), .A2(B[5]), .ZN(n444) );
  NAND2_X1 U558 ( .A1(A[5]), .A2(B[5]), .ZN(n79) );
  NAND2_X1 U559 ( .A1(n307), .A2(n294), .ZN(n306) );
  NAND4_X1 U560 ( .A1(net507278), .A2(net507279), .A3(net507280), .A4(n29), 
        .ZN(net537591) );
  NAND4_X1 U561 ( .A1(net507278), .A2(net507279), .A3(net507280), .A4(n29), 
        .ZN(net507122) );
  NAND4_X1 U562 ( .A1(n407), .A2(n411), .A3(n419), .A4(n57), .ZN(n383) );
  INV_X1 U563 ( .A(n383), .ZN(n506) );
  AOI21_X1 U564 ( .B1(n381), .B2(n382), .A(n383), .ZN(n378) );
  NOR2_X1 U565 ( .A1(n199), .A2(n200), .ZN(n198) );
  OAI221_X1 U566 ( .B1(n543), .B2(n297), .C1(n490), .C2(n200), .A(n298), .ZN(
        n20) );
  NAND2_X1 U568 ( .A1(n298), .A2(n295), .ZN(n305) );
  OAI221_X1 U569 ( .B1(n543), .B2(n297), .C1(n490), .C2(n200), .A(n298), .ZN(
        n272) );
  NAND2_X1 U570 ( .A1(n294), .A2(n295), .ZN(n297) );
  NAND4_X1 U571 ( .A1(n292), .A2(n293), .A3(n294), .A4(n295), .ZN(n200) );
  NOR2_X1 U572 ( .A1(n201), .A2(n465), .ZN(n197) );
  INV_X1 U573 ( .A(n465), .ZN(n536) );
  NAND2_X1 U575 ( .A1(n247), .A2(n248), .ZN(n258) );
  OAI21_X1 U576 ( .B1(n489), .B2(n202), .A(n221), .ZN(n247) );
  INV_X1 U577 ( .A(n26), .ZN(n501) );
  OAI21_X1 U580 ( .B1(n468), .B2(n544), .A(n302), .ZN(n307) );
  XNOR2_X1 U581 ( .A(n304), .B(n305), .ZN(SUM[35]) );
  NAND2_X1 U582 ( .A1(n303), .A2(n306), .ZN(n304) );
  NAND2_X1 U584 ( .A1(n466), .A2(n454), .ZN(n235) );
  NAND2_X1 U586 ( .A1(n209), .A2(n227), .ZN(n226) );
  NAND2_X1 U587 ( .A1(n272), .A2(n271), .ZN(n290) );
  XNOR2_X1 U588 ( .A(n253), .B(n472), .ZN(SUM[42]) );
  NAND2_X1 U589 ( .A1(n243), .A2(n252), .ZN(n251) );
endmodule


module RCA_NBIT64_14 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_14_DW01_add_6 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), 
        .SUM({Co, S}) );
endmodule


module RCA_NBIT64_13_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net497441, net497398, net497394, net497392, net497381, net497376,
         net497375, net497373, net497366, net497362, net497361, net497359,
         net497352, net497349, net497348, net497347, net497338, net497337,
         net497317, net497316, net497312, net497311, net497310, net497309,
         net497287, net497282, net497280, net497278, net497268, net497267,
         net497262, net497254, net497253, net497252, net497251, net497240,
         net497239, net497238, net497236, net497232, net497231, net497222,
         net497212, net497205, net497196, net497195, net497194, net497193,
         net497192, net497189, net497188, net497187, net497156, net497148,
         net497147, net497146, net497143, net497070, net497069, net497068,
         net497062, net534733, net535589, net537101, net537534, net537813,
         net538090, net538199, net538264, net538609, net538905, net497165,
         net497190, net497186, net497078, net497066, net537617, net497390,
         net497224, net537913, net497245, net497234, net497233, net497225,
         net497219, net497218, net497217, net497216, net497197, net537151,
         net535368, net497250, net497249, net497244, net497243, net497166,
         net497149, net497167, net497155, net497154, net497153, net497152,
         net497151, n1, n2, n4, n5, n8, n9, n10, n11, n12, n13, n14, n17, n18,
         n21, n23, n24, n26, n27, n29, n31, n33, n34, n36, n39, n41, n42, n44,
         n47, n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n75, n76, n77,
         n78, n80, n81, n82, n83, n84, n85, n88, n89, n92, n93, n95, n96, n97,
         n99, n100, n101, n102, n103, n104, n105, n107, n108, n109, n111, n112,
         n113, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n129, n131, n132, n134, n135, n136, n138, n139, n140,
         n142, n143, n144, n147, n148, n149, n150, n151, n152, n153, n157,
         n158, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n174, n176, n177, n178, n179, n180, n181, n182,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n198, n199, n200, n201, n202, n203, n205, n206, n207, n209,
         n210, n211, n212, n214, n216, n217, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n237, n239, n240, n241, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n259, n260, n261, n262,
         n263, n264, n265, n266, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n295, n296, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n314,
         n315, n316, n317, n318, n319, n320, n322, n323, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n360, n361,
         n362, n363, n364, n365, n366, n368, n369, n372, n373, n375, n376,
         n377, n378, n379, n381, n382, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n394, n395, n396, n397, n398, n399, n400, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513;

  OR2_X2 U8 ( .A1(B[14]), .A2(A[14]), .ZN(n351) );
  NAND3_X1 U11 ( .A1(net497282), .A2(net538905), .A3(n5), .ZN(net497280) );
  NAND3_X1 U13 ( .A1(net497231), .A2(n417), .A3(n9), .ZN(net497390) );
  OR2_X2 U15 ( .A1(B[42]), .A2(A[42]), .ZN(n226) );
  OR2_X2 U34 ( .A1(A[22]), .A2(B[22]), .ZN(net497348) );
  OR2_X2 U35 ( .A1(B[38]), .A2(A[38]), .ZN(net497153) );
  NAND3_X1 U44 ( .A1(net497348), .A2(net497349), .A3(net497338), .ZN(n273) );
  XOR2_X1 U49 ( .A(net538090), .B(n250), .Z(SUM[33]) );
  NAND3_X1 U95 ( .A1(net497287), .A2(net497254), .A3(net497249), .ZN(net538609) );
  NAND3_X1 U101 ( .A1(net497218), .A2(net497216), .A3(net497217), .ZN(
        net497197) );
  NAND3_X1 U118 ( .A1(net497347), .A2(n483), .A3(n502), .ZN(n33) );
  NAND3_X1 U127 ( .A1(net534733), .A2(net497398), .A3(n484), .ZN(net497394) );
  OR2_X2 U155 ( .A1(A[26]), .A2(B[26]), .ZN(net497253) );
  OR2_X2 U156 ( .A1(A[23]), .A2(B[23]), .ZN(net497349) );
  NAND3_X1 U160 ( .A1(n352), .A2(n351), .A3(n4), .ZN(n350) );
  OR2_X2 U161 ( .A1(B[12]), .A2(A[12]), .ZN(n335) );
  OR2_X2 U162 ( .A1(A[13]), .A2(B[13]), .ZN(n334) );
  NOR2_X2 U166 ( .A1(A[16]), .A2(B[16]), .ZN(net537101) );
  OR2_X2 U172 ( .A1(A[19]), .A2(B[19]), .ZN(net497231) );
  OR2_X2 U349 ( .A1(B[20]), .A2(A[20]), .ZN(net497347) );
  NAND3_X1 U440 ( .A1(n317), .A2(net538199), .A3(n318), .ZN(n316) );
  NAND3_X1 U530 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n163) );
  NAND3_X1 U554 ( .A1(net497252), .A2(n279), .A3(net497253), .ZN(n263) );
  NAND3_X1 U555 ( .A1(net497254), .A2(net538905), .A3(n49), .ZN(n261) );
  NAND3_X1 U562 ( .A1(n290), .A2(n289), .A3(n483), .ZN(net497311) );
  NAND3_X1 U574 ( .A1(net497232), .A2(net497347), .A3(net497231), .ZN(n296) );
  NAND3_X1 U576 ( .A1(n409), .A2(B[17]), .A3(net497398), .ZN(n304) );
  NAND3_X1 U582 ( .A1(n44), .A2(n340), .A3(n58), .ZN(n343) );
  NAND3_X1 U583 ( .A1(n344), .A2(n345), .A3(n246), .ZN(n341) );
  NAND3_X1 U584 ( .A1(n349), .A2(n346), .A3(n350), .ZN(n348) );
  NAND3_X1 U585 ( .A1(n351), .A2(n353), .A3(n334), .ZN(n349) );
  NAND3_X1 U589 ( .A1(n361), .A2(n366), .A3(n338), .ZN(n352) );
  NAND3_X1 U590 ( .A1(n369), .A2(n61), .A3(n368), .ZN(n366) );
  NAND3_X1 U596 ( .A1(n385), .A2(n386), .A3(n384), .ZN(n382) );
  NAND3_X1 U601 ( .A1(n385), .A2(n63), .A3(n386), .ZN(n57) );
  NAND3_X1 U602 ( .A1(n62), .A2(n71), .A3(n373), .ZN(n386) );
  NAND3_X1 U603 ( .A1(n392), .A2(n391), .A3(n390), .ZN(n373) );
  NAND3_X1 U604 ( .A1(n76), .A2(n509), .A3(n68), .ZN(n391) );
  NAND3_X1 U606 ( .A1(n44), .A2(n123), .A3(n345), .ZN(n385) );
  OR2_X2 U6 ( .A1(B[27]), .A2(A[27]), .ZN(net497254) );
  AND2_X2 U22 ( .A1(n484), .A2(n487), .ZN(n9) );
  OR2_X2 U76 ( .A1(B[37]), .A2(A[37]), .ZN(net497151) );
  OR2_X2 U173 ( .A1(B[25]), .A2(A[25]), .ZN(net497252) );
  AND2_X2 U352 ( .A1(B[16]), .A2(A[16]), .ZN(net534733) );
  OR2_X2 U390 ( .A1(B[34]), .A2(A[34]), .ZN(net497188) );
  CLKBUF_X1 U2 ( .A(A[7]), .Z(n403) );
  NAND2_X1 U3 ( .A1(B[20]), .A2(A[20]), .ZN(n286) );
  INV_X1 U4 ( .A(net537101), .ZN(n487) );
  OR2_X1 U5 ( .A1(B[24]), .A2(A[24]), .ZN(net497251) );
  OR2_X1 U7 ( .A1(B[28]), .A2(A[28]), .ZN(net497249) );
  AND2_X1 U9 ( .A1(net497212), .A2(net497192), .ZN(net538090) );
  AND2_X1 U10 ( .A1(n400), .A2(n397), .ZN(SUM[0]) );
  OR2_X1 U12 ( .A1(B[29]), .A2(A[29]), .ZN(net497250) );
  OR2_X1 U14 ( .A1(B[40]), .A2(A[40]), .ZN(n229) );
  OR2_X1 U16 ( .A1(B[41]), .A2(A[41]), .ZN(n225) );
  OR2_X1 U17 ( .A1(B[39]), .A2(A[39]), .ZN(net497147) );
  OR2_X1 U18 ( .A1(B[36]), .A2(A[36]), .ZN(net497156) );
  OR2_X1 U19 ( .A1(B[32]), .A2(A[32]), .ZN(net497195) );
  OR2_X1 U20 ( .A1(B[44]), .A2(A[44]), .ZN(n198) );
  OR2_X1 U21 ( .A1(B[46]), .A2(A[46]), .ZN(n200) );
  OR2_X1 U23 ( .A1(B[50]), .A2(A[50]), .ZN(n170) );
  OR2_X1 U24 ( .A1(B[49]), .A2(A[49]), .ZN(n168) );
  OR2_X1 U25 ( .A1(B[48]), .A2(A[48]), .ZN(n167) );
  OR2_X1 U26 ( .A1(B[52]), .A2(A[52]), .ZN(n149) );
  OR2_X1 U27 ( .A1(B[55]), .A2(A[55]), .ZN(n148) );
  OR2_X1 U28 ( .A1(B[54]), .A2(A[54]), .ZN(n147) );
  OR2_X1 U29 ( .A1(B[53]), .A2(A[53]), .ZN(n150) );
  OR2_X1 U30 ( .A1(B[56]), .A2(A[56]), .ZN(n118) );
  OR2_X1 U31 ( .A1(B[58]), .A2(A[58]), .ZN(n116) );
  OR2_X1 U32 ( .A1(B[57]), .A2(A[57]), .ZN(n119) );
  OR2_X1 U33 ( .A1(A[9]), .A2(B[9]), .ZN(n58) );
  AND3_X1 U36 ( .A1(n495), .A2(net497245), .A3(n483), .ZN(n404) );
  AND3_X1 U37 ( .A1(n457), .A2(net497070), .A3(n462), .ZN(n405) );
  AND2_X1 U38 ( .A1(n225), .A2(n229), .ZN(n406) );
  CLKBUF_X1 U39 ( .A(net535589), .Z(n407) );
  CLKBUF_X1 U40 ( .A(net497197), .Z(n408) );
  CLKBUF_X1 U41 ( .A(A[17]), .Z(n409) );
  OR2_X1 U42 ( .A1(B[8]), .A2(A[8]), .ZN(n44) );
  OR2_X1 U43 ( .A1(A[15]), .A2(B[15]), .ZN(n410) );
  OR2_X1 U45 ( .A1(A[15]), .A2(B[15]), .ZN(n336) );
  AND3_X2 U46 ( .A1(n319), .A2(n317), .A3(n318), .ZN(net535589) );
  AND3_X1 U47 ( .A1(net497349), .A2(net497348), .A3(n8), .ZN(net537617) );
  CLKBUF_X1 U48 ( .A(n59), .Z(n411) );
  NAND2_X1 U50 ( .A1(net535368), .A2(n404), .ZN(net497216) );
  OR2_X1 U51 ( .A1(A[35]), .A2(B[35]), .ZN(net497189) );
  NAND4_X1 U52 ( .A1(n304), .A2(net497394), .A3(n305), .A4(n306), .ZN(n412) );
  OR2_X1 U53 ( .A1(A[31]), .A2(B[31]), .ZN(n413) );
  AND2_X1 U54 ( .A1(n216), .A2(n205), .ZN(n414) );
  NAND2_X1 U55 ( .A1(net537617), .A2(n481), .ZN(n415) );
  NAND2_X1 U56 ( .A1(n51), .A2(n405), .ZN(n192) );
  CLKBUF_X1 U57 ( .A(n70), .Z(n416) );
  NOR2_X1 U58 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  OR2_X1 U59 ( .A1(B[18]), .A2(A[18]), .ZN(n417) );
  OR2_X1 U60 ( .A1(A[18]), .A2(B[18]), .ZN(net497398) );
  OR2_X1 U61 ( .A1(A[33]), .A2(B[33]), .ZN(net497196) );
  NAND3_X1 U62 ( .A1(n221), .A2(n226), .A3(n406), .ZN(n195) );
  OR2_X1 U63 ( .A1(A[43]), .A2(B[43]), .ZN(n221) );
  NAND2_X1 U64 ( .A1(n483), .A2(net497381), .ZN(n34) );
  XNOR2_X1 U65 ( .A(n18), .B(n418), .ZN(SUM[35]) );
  NAND2_X1 U66 ( .A1(net497187), .A2(net497189), .ZN(n418) );
  XNOR2_X1 U67 ( .A(n268), .B(n419), .ZN(SUM[27]) );
  NAND2_X1 U68 ( .A1(net497254), .A2(n274), .ZN(n419) );
  AND4_X1 U69 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n51) );
  XNOR2_X1 U70 ( .A(n420), .B(net537813), .ZN(SUM[38]) );
  NAND2_X1 U71 ( .A1(net497153), .A2(net497149), .ZN(n420) );
  AND2_X1 U72 ( .A1(n216), .A2(n205), .ZN(n421) );
  XOR2_X1 U73 ( .A(n23), .B(n320), .Z(SUM[17]) );
  XNOR2_X1 U74 ( .A(n408), .B(n422), .ZN(SUM[32]) );
  NAND2_X1 U75 ( .A1(net497192), .A2(net497195), .ZN(n422) );
  XOR2_X1 U77 ( .A(n352), .B(n423), .Z(SUM[12]) );
  AND2_X1 U78 ( .A1(n325), .A2(n335), .ZN(n423) );
  XOR2_X1 U79 ( .A(n424), .B(n153), .Z(SUM[54]) );
  AND2_X1 U80 ( .A1(n147), .A2(n144), .ZN(n424) );
  XOR2_X1 U81 ( .A(n425), .B(n182), .Z(SUM[50]) );
  AND2_X1 U82 ( .A1(n170), .A2(n177), .ZN(n425) );
  XOR2_X1 U83 ( .A(n260), .B(n426), .Z(SUM[28]) );
  AND2_X1 U84 ( .A1(net497249), .A2(net497238), .ZN(n426) );
  XOR2_X1 U85 ( .A(net538264), .B(n427), .Z(SUM[36]) );
  AND2_X1 U86 ( .A1(net497156), .A2(net497155), .ZN(n427) );
  XNOR2_X1 U87 ( .A(n428), .B(n209), .ZN(SUM[47]) );
  NAND2_X1 U88 ( .A1(n191), .A2(n201), .ZN(n428) );
  XOR2_X1 U89 ( .A(n429), .B(n251), .Z(SUM[31]) );
  AND2_X1 U90 ( .A1(n413), .A2(net497236), .ZN(n429) );
  NAND2_X1 U91 ( .A1(n482), .A2(n502), .ZN(net497361) );
  AOI21_X1 U92 ( .B1(net497066), .B2(n450), .A(n449), .ZN(net497062) );
  INV_X1 U93 ( .A(net497068), .ZN(n449) );
  INV_X1 U94 ( .A(net497390), .ZN(n483) );
  OAI21_X1 U96 ( .B1(n493), .B2(net497219), .A(net535368), .ZN(net497218) );
  AOI21_X1 U97 ( .B1(net497233), .B2(net497234), .A(n498), .ZN(net497217) );
  INV_X1 U98 ( .A(n134), .ZN(n437) );
  INV_X1 U99 ( .A(n296), .ZN(n482) );
  NOR2_X1 U100 ( .A1(n407), .A2(n491), .ZN(net497245) );
  INV_X1 U102 ( .A(A[11]), .ZN(n448) );
  INV_X1 U103 ( .A(n103), .ZN(n436) );
  INV_X1 U104 ( .A(net497366), .ZN(n502) );
  INV_X1 U105 ( .A(net497078), .ZN(n462) );
  NAND2_X1 U106 ( .A1(n482), .A2(n289), .ZN(net497376) );
  INV_X1 U107 ( .A(net497224), .ZN(n495) );
  INV_X1 U108 ( .A(net497352), .ZN(n481) );
  INV_X1 U109 ( .A(net497222), .ZN(n493) );
  INV_X1 U110 ( .A(net497309), .ZN(n496) );
  INV_X1 U111 ( .A(n271), .ZN(n497) );
  NOR2_X1 U112 ( .A1(n78), .A2(n469), .ZN(SUM[64]) );
  AND2_X1 U113 ( .A1(n417), .A2(n306), .ZN(n10) );
  NAND4_X1 U114 ( .A1(n148), .A2(n147), .A3(n149), .A4(n150), .ZN(n136) );
  AOI21_X1 U115 ( .B1(n139), .B2(n140), .A(n54), .ZN(n138) );
  OAI211_X1 U116 ( .C1(n477), .C2(n142), .A(n143), .B(n144), .ZN(n140) );
  NAND2_X1 U117 ( .A1(net497251), .A2(n265), .ZN(n283) );
  NAND2_X1 U119 ( .A1(net497250), .A2(net497239), .ZN(net497278) );
  NAND2_X1 U120 ( .A1(n289), .A2(n287), .ZN(n300) );
  NAND2_X1 U121 ( .A1(net497347), .A2(n483), .ZN(n302) );
  NAND2_X1 U122 ( .A1(n150), .A2(n143), .ZN(n158) );
  XOR2_X1 U123 ( .A(n430), .B(n217), .Z(SUM[44]) );
  AND2_X1 U124 ( .A1(n198), .A2(n205), .ZN(n430) );
  NAND2_X1 U125 ( .A1(n200), .A2(n207), .ZN(n212) );
  NAND2_X1 U126 ( .A1(n149), .A2(n142), .ZN(n161) );
  NAND2_X1 U128 ( .A1(n226), .A2(n223), .ZN(n234) );
  NOR2_X1 U129 ( .A1(n451), .A2(n452), .ZN(n26) );
  INV_X1 U130 ( .A(net497154), .ZN(n451) );
  NOR2_X1 U131 ( .A1(n492), .A2(n494), .ZN(n276) );
  INV_X1 U132 ( .A(n266), .ZN(n492) );
  OAI21_X1 U133 ( .B1(n252), .B2(net497262), .A(net497240), .ZN(n251) );
  NAND2_X1 U134 ( .A1(net497231), .A2(n305), .ZN(n308) );
  NAND2_X1 U135 ( .A1(n417), .A2(n9), .ZN(n310) );
  OAI211_X1 U136 ( .C1(n34), .C2(net535589), .A(net497375), .B(net497376), 
        .ZN(net497373) );
  AOI21_X1 U137 ( .B1(n490), .B2(n289), .A(n504), .ZN(net497375) );
  INV_X1 U138 ( .A(net534733), .ZN(n486) );
  INV_X1 U139 ( .A(n149), .ZN(n478) );
  NAND2_X1 U140 ( .A1(net497196), .A2(net497193), .ZN(n250) );
  INV_X1 U141 ( .A(n225), .ZN(n458) );
  OAI21_X1 U142 ( .B1(n432), .B2(n477), .A(n143), .ZN(n153) );
  OAI21_X1 U143 ( .B1(n433), .B2(n468), .A(n112), .ZN(n127) );
  INV_X1 U144 ( .A(n131), .ZN(n433) );
  OAI21_X1 U145 ( .B1(n436), .B2(n472), .A(n89), .ZN(n100) );
  OAI21_X1 U146 ( .B1(n435), .B2(n471), .A(n88), .ZN(n96) );
  INV_X1 U147 ( .A(n100), .ZN(n435) );
  OAI21_X1 U148 ( .B1(n473), .B2(n437), .A(n111), .ZN(n131) );
  INV_X1 U149 ( .A(n118), .ZN(n473) );
  NAND2_X1 U150 ( .A1(n44), .A2(n63), .ZN(n60) );
  NOR2_X1 U151 ( .A1(net534733), .A2(net537101), .ZN(n328) );
  NAND2_X1 U152 ( .A1(n340), .A2(n377), .ZN(n387) );
  NAND2_X1 U153 ( .A1(net497349), .A2(net497316), .ZN(n291) );
  OAI211_X1 U154 ( .C1(n33), .C2(net535589), .A(net497361), .B(net497362), 
        .ZN(net497359) );
  INV_X1 U157 ( .A(n314), .ZN(n485) );
  NAND2_X1 U158 ( .A1(n222), .A2(n223), .ZN(n220) );
  NOR2_X1 U159 ( .A1(n12), .A2(n224), .ZN(n219) );
  AND2_X1 U163 ( .A1(n227), .A2(n228), .ZN(n12) );
  OAI21_X1 U164 ( .B1(n431), .B2(n464), .A(n178), .ZN(n182) );
  OAI211_X1 U165 ( .C1(n506), .C2(n325), .A(n326), .B(n346), .ZN(n323) );
  NAND4_X1 U167 ( .A1(n190), .A2(n191), .A3(n192), .A4(n193), .ZN(n166) );
  NAND2_X1 U168 ( .A1(n202), .A2(n203), .ZN(n190) );
  NAND2_X1 U169 ( .A1(n51), .A2(n194), .ZN(n193) );
  XNOR2_X1 U170 ( .A(n135), .B(n134), .ZN(SUM[56]) );
  NAND2_X1 U171 ( .A1(n118), .A2(n111), .ZN(n135) );
  AND2_X1 U174 ( .A1(n36), .A2(net497347), .ZN(n8) );
  XNOR2_X1 U175 ( .A(n187), .B(n185), .ZN(SUM[49]) );
  NAND2_X1 U176 ( .A1(n168), .A2(n178), .ZN(n187) );
  XNOR2_X1 U177 ( .A(n237), .B(n440), .ZN(SUM[41]) );
  NAND2_X1 U178 ( .A1(n225), .A2(n227), .ZN(n237) );
  XNOR2_X1 U179 ( .A(n303), .B(net497392), .ZN(SUM[20]) );
  NAND2_X1 U180 ( .A1(net497347), .A2(n286), .ZN(n303) );
  OAI21_X1 U181 ( .B1(net535589), .B2(net497390), .A(net497352), .ZN(net497392) );
  XNOR2_X1 U182 ( .A(n179), .B(n180), .ZN(SUM[51]) );
  NAND2_X1 U183 ( .A1(n169), .A2(n174), .ZN(n179) );
  XNOR2_X1 U184 ( .A(n132), .B(n131), .ZN(SUM[57]) );
  NAND2_X1 U185 ( .A1(n119), .A2(n112), .ZN(n132) );
  XNOR2_X1 U186 ( .A(n129), .B(n127), .ZN(SUM[58]) );
  NAND2_X1 U187 ( .A1(n116), .A2(n113), .ZN(n129) );
  XNOR2_X1 U188 ( .A(n104), .B(n103), .ZN(SUM[60]) );
  NAND2_X1 U189 ( .A1(n102), .A2(n89), .ZN(n104) );
  XNOR2_X1 U190 ( .A(n101), .B(n100), .ZN(SUM[61]) );
  NAND2_X1 U191 ( .A1(n99), .A2(n88), .ZN(n101) );
  XNOR2_X1 U192 ( .A(n97), .B(n96), .ZN(SUM[62]) );
  NAND2_X1 U193 ( .A1(n95), .A2(n85), .ZN(n97) );
  NAND2_X1 U194 ( .A1(n261), .A2(net497222), .ZN(n260) );
  XNOR2_X1 U195 ( .A(n414), .B(n214), .ZN(SUM[45]) );
  NOR2_X1 U196 ( .A1(n453), .A2(n454), .ZN(n214) );
  INV_X1 U197 ( .A(n206), .ZN(n453) );
  XNOR2_X1 U198 ( .A(n439), .B(n239), .ZN(SUM[40]) );
  NOR2_X1 U199 ( .A1(n455), .A2(n456), .ZN(n239) );
  INV_X1 U200 ( .A(n229), .ZN(n456) );
  XNOR2_X1 U201 ( .A(n125), .B(n126), .ZN(SUM[59]) );
  NOR2_X1 U202 ( .A1(n465), .A2(n55), .ZN(n126) );
  AOI21_X1 U203 ( .B1(n116), .B2(n127), .A(n467), .ZN(n125) );
  INV_X1 U204 ( .A(n113), .ZN(n467) );
  NAND4_X1 U205 ( .A1(net497251), .A2(net497252), .A3(net497253), .A4(
        net497254), .ZN(net497224) );
  NAND4_X1 U206 ( .A1(net497195), .A2(net497196), .A3(net497188), .A4(
        net497189), .ZN(net497078) );
  OAI21_X1 U207 ( .B1(n461), .B2(net497186), .A(net497187), .ZN(net497066) );
  XNOR2_X1 U208 ( .A(n92), .B(n93), .ZN(SUM[63]) );
  NAND2_X1 U209 ( .A1(n84), .A2(n80), .ZN(n92) );
  OAI21_X1 U210 ( .B1(n434), .B2(n470), .A(n85), .ZN(n93) );
  INV_X1 U211 ( .A(n96), .ZN(n434) );
  OAI211_X1 U212 ( .C1(n464), .C2(n176), .A(n177), .B(n178), .ZN(n172) );
  OAI211_X1 U213 ( .C1(n499), .C2(net497238), .A(net497239), .B(net497240), 
        .ZN(net497234) );
  OAI211_X1 U214 ( .C1(n454), .C2(n205), .A(n206), .B(n207), .ZN(n203) );
  OAI21_X1 U215 ( .B1(n421), .B2(n454), .A(n206), .ZN(n211) );
  OAI21_X1 U216 ( .B1(n444), .B2(n269), .A(n266), .ZN(n268) );
  XNOR2_X1 U217 ( .A(n354), .B(n355), .ZN(SUM[14]) );
  NAND2_X1 U218 ( .A1(n351), .A2(n346), .ZN(n354) );
  OAI21_X1 U219 ( .B1(n39), .B2(n357), .A(n358), .ZN(n356) );
  XNOR2_X1 U220 ( .A(n281), .B(n280), .ZN(SUM[25]) );
  NAND2_X1 U221 ( .A1(net497252), .A2(n264), .ZN(n280) );
  OAI211_X1 U222 ( .C1(net537101), .C2(net538199), .A(net497441), .B(n13), 
        .ZN(n23) );
  OR2_X1 U223 ( .A1(net537101), .A2(n318), .ZN(n13) );
  OAI21_X1 U224 ( .B1(n105), .B2(n437), .A(n107), .ZN(n103) );
  NAND4_X1 U225 ( .A1(n117), .A2(n116), .A3(n118), .A4(n119), .ZN(n105) );
  AOI21_X1 U226 ( .B1(n108), .B2(n109), .A(n55), .ZN(n107) );
  OAI211_X1 U227 ( .C1(n468), .C2(n111), .A(n112), .B(n113), .ZN(n109) );
  XNOR2_X1 U228 ( .A(n189), .B(n166), .ZN(SUM[48]) );
  NAND2_X1 U229 ( .A1(n167), .A2(n176), .ZN(n189) );
  NAND2_X1 U230 ( .A1(n510), .A2(n503), .ZN(n289) );
  XNOR2_X1 U231 ( .A(net497166), .B(net497165), .ZN(SUM[39]) );
  NAND2_X1 U232 ( .A1(net497148), .A2(net497147), .ZN(net497165) );
  NAND2_X1 U233 ( .A1(net497167), .A2(net497149), .ZN(net497166) );
  XNOR2_X1 U234 ( .A(n231), .B(n230), .ZN(SUM[43]) );
  XNOR2_X1 U235 ( .A(n151), .B(n152), .ZN(SUM[55]) );
  NOR2_X1 U236 ( .A1(n474), .A2(n54), .ZN(n152) );
  AOI21_X1 U237 ( .B1(n147), .B2(n153), .A(n476), .ZN(n151) );
  INV_X1 U238 ( .A(n144), .ZN(n476) );
  NOR2_X1 U239 ( .A1(n446), .A2(n52), .ZN(n379) );
  AOI21_X1 U240 ( .B1(n381), .B2(n382), .A(n447), .ZN(n378) );
  INV_X1 U241 ( .A(n338), .ZN(n446) );
  NAND2_X1 U242 ( .A1(n345), .A2(n123), .ZN(n372) );
  AOI21_X1 U243 ( .B1(n312), .B2(n417), .A(n489), .ZN(n311) );
  INV_X1 U244 ( .A(n306), .ZN(n489) );
  INV_X1 U245 ( .A(net497156), .ZN(n459) );
  XNOR2_X1 U246 ( .A(n348), .B(n347), .ZN(SUM[15]) );
  NOR2_X1 U247 ( .A1(n31), .A2(net497224), .ZN(net497219) );
  NOR2_X1 U248 ( .A1(n480), .A2(n488), .ZN(net497225) );
  INV_X1 U249 ( .A(net497316), .ZN(n500) );
  AOI21_X1 U250 ( .B1(n171), .B2(n172), .A(n463), .ZN(n162) );
  AND2_X1 U251 ( .A1(n167), .A2(n168), .ZN(n165) );
  NOR2_X1 U252 ( .A1(n292), .A2(n293), .ZN(net497362) );
  OAI21_X1 U253 ( .B1(n501), .B2(n287), .A(n288), .ZN(n293) );
  NOR2_X1 U254 ( .A1(n286), .A2(net497366), .ZN(n292) );
  NAND2_X1 U255 ( .A1(n279), .A2(net497252), .ZN(net497309) );
  NAND2_X1 U256 ( .A1(net497231), .A2(n412), .ZN(net497352) );
  NOR2_X1 U257 ( .A1(n506), .A2(n505), .ZN(n358) );
  INV_X1 U258 ( .A(n335), .ZN(n505) );
  NOR2_X1 U259 ( .A1(n376), .A2(n48), .ZN(n381) );
  NOR2_X1 U260 ( .A1(n474), .A2(n475), .ZN(n139) );
  INV_X1 U261 ( .A(n147), .ZN(n475) );
  NOR2_X1 U262 ( .A1(n465), .A2(n466), .ZN(n108) );
  INV_X1 U263 ( .A(n116), .ZN(n466) );
  NOR2_X1 U264 ( .A1(n48), .A2(n53), .ZN(n369) );
  INV_X1 U265 ( .A(n199), .ZN(n454) );
  XNOR2_X1 U266 ( .A(n363), .B(n362), .ZN(SUM[13]) );
  NAND2_X1 U267 ( .A1(n334), .A2(n326), .ZN(n362) );
  OAI21_X1 U268 ( .B1(n39), .B2(n365), .A(n335), .ZN(n364) );
  NAND2_X1 U269 ( .A1(n510), .A2(n503), .ZN(n36) );
  NAND2_X1 U270 ( .A1(net497287), .A2(net497254), .ZN(net497222) );
  NAND2_X1 U271 ( .A1(net497251), .A2(net497252), .ZN(n271) );
  NAND2_X1 U272 ( .A1(n337), .A2(n338), .ZN(n330) );
  NAND2_X1 U273 ( .A1(n47), .A2(n323), .ZN(n317) );
  AND2_X1 U274 ( .A1(n445), .A2(n448), .ZN(n53) );
  OAI211_X1 U275 ( .C1(n329), .C2(n330), .A(n2), .B(n332), .ZN(net538199) );
  NAND2_X1 U276 ( .A1(n262), .A2(n263), .ZN(net497287) );
  AND2_X1 U277 ( .A1(n274), .A2(n266), .ZN(n262) );
  NAND2_X1 U278 ( .A1(n264), .A2(n265), .ZN(n279) );
  INV_X1 U279 ( .A(net497151), .ZN(n452) );
  INV_X1 U280 ( .A(n287), .ZN(n504) );
  NAND2_X1 U281 ( .A1(n360), .A2(n361), .ZN(n357) );
  AND2_X1 U282 ( .A1(n325), .A2(n338), .ZN(n360) );
  INV_X1 U283 ( .A(n99), .ZN(n471) );
  INV_X1 U284 ( .A(n95), .ZN(n470) );
  INV_X1 U285 ( .A(n148), .ZN(n474) );
  INV_X1 U286 ( .A(n117), .ZN(n465) );
  INV_X1 U287 ( .A(n102), .ZN(n472) );
  NAND2_X1 U288 ( .A1(n361), .A2(n338), .ZN(n365) );
  INV_X1 U289 ( .A(n150), .ZN(n477) );
  INV_X1 U290 ( .A(n119), .ZN(n468) );
  INV_X1 U291 ( .A(n334), .ZN(n506) );
  INV_X1 U292 ( .A(n168), .ZN(n464) );
  INV_X1 U293 ( .A(net497232), .ZN(n480) );
  AND3_X1 U294 ( .A1(net497252), .A2(net497251), .A3(net497253), .ZN(net538905) );
  AND2_X1 U295 ( .A1(n445), .A2(n448), .ZN(n52) );
  AND2_X1 U296 ( .A1(n413), .A2(net537151), .ZN(net535368) );
  AND2_X1 U297 ( .A1(net538609), .A2(net497238), .ZN(n41) );
  NAND2_X1 U298 ( .A1(n270), .A2(net497253), .ZN(n269) );
  NAND2_X1 U299 ( .A1(n271), .A2(net497309), .ZN(n270) );
  INV_X1 U300 ( .A(net497196), .ZN(n479) );
  NAND2_X1 U301 ( .A1(n225), .A2(n226), .ZN(n224) );
  AND2_X1 U302 ( .A1(n334), .A2(n335), .ZN(n4) );
  INV_X1 U303 ( .A(n228), .ZN(n455) );
  INV_X1 U304 ( .A(net497250), .ZN(n499) );
  NAND2_X1 U305 ( .A1(n326), .A2(n325), .ZN(n353) );
  INV_X1 U306 ( .A(n286), .ZN(n490) );
  INV_X1 U307 ( .A(net497236), .ZN(n498) );
  AND2_X1 U308 ( .A1(n273), .A2(net497316), .ZN(n284) );
  AND2_X1 U309 ( .A1(net497347), .A2(n36), .ZN(net497381) );
  INV_X1 U310 ( .A(n174), .ZN(n463) );
  AND3_X1 U311 ( .A1(net497151), .A2(net497152), .A3(net497153), .ZN(n11) );
  NAND2_X1 U312 ( .A1(net497148), .A2(net497149), .ZN(net497146) );
  NAND2_X1 U313 ( .A1(net497154), .A2(net497155), .ZN(net497152) );
  INV_X1 U314 ( .A(net497253), .ZN(n494) );
  INV_X1 U315 ( .A(net497231), .ZN(n488) );
  AND2_X1 U316 ( .A1(n170), .A2(n169), .ZN(n171) );
  INV_X1 U317 ( .A(n377), .ZN(n447) );
  AND2_X1 U318 ( .A1(net497254), .A2(net497249), .ZN(n5) );
  AND2_X1 U319 ( .A1(net497337), .A2(net497338), .ZN(net537913) );
  AND2_X1 U320 ( .A1(n41), .A2(n42), .ZN(n252) );
  AND2_X1 U321 ( .A1(net497239), .A2(net497280), .ZN(n42) );
  NAND2_X1 U322 ( .A1(n394), .A2(n68), .ZN(n390) );
  AND2_X1 U323 ( .A1(n70), .A2(n66), .ZN(n392) );
  AND2_X1 U324 ( .A1(n169), .A2(n170), .ZN(n164) );
  XNOR2_X1 U325 ( .A(n64), .B(n65), .ZN(SUM[7]) );
  NAND2_X1 U326 ( .A1(n66), .A2(n67), .ZN(n65) );
  NAND2_X1 U327 ( .A1(n416), .A2(n71), .ZN(n64) );
  NAND2_X1 U328 ( .A1(n68), .A2(n69), .ZN(n67) );
  XNOR2_X1 U329 ( .A(n186), .B(n123), .ZN(SUM[4]) );
  NAND2_X1 U330 ( .A1(n122), .A2(n124), .ZN(n186) );
  XNOR2_X1 U331 ( .A(n240), .B(n241), .ZN(SUM[3]) );
  OAI21_X1 U332 ( .B1(n512), .B2(n511), .A(n244), .ZN(n241) );
  NAND2_X1 U333 ( .A1(n246), .A2(n247), .ZN(n240) );
  INV_X1 U334 ( .A(n245), .ZN(n512) );
  XNOR2_X1 U335 ( .A(n254), .B(n245), .ZN(SUM[2]) );
  NAND2_X1 U336 ( .A1(n259), .A2(n244), .ZN(n254) );
  XNOR2_X1 U337 ( .A(n72), .B(n69), .ZN(SUM[6]) );
  NAND2_X1 U338 ( .A1(n68), .A2(n66), .ZN(n72) );
  XNOR2_X1 U339 ( .A(n120), .B(n77), .ZN(SUM[5]) );
  NAND2_X1 U340 ( .A1(n76), .A2(n75), .ZN(n120) );
  XNOR2_X1 U341 ( .A(n307), .B(n513), .ZN(SUM[1]) );
  NAND2_X1 U342 ( .A1(n257), .A2(n256), .ZN(n307) );
  OAI21_X1 U343 ( .B1(n508), .B2(n507), .A(n75), .ZN(n69) );
  INV_X1 U344 ( .A(n77), .ZN(n508) );
  INV_X1 U345 ( .A(n76), .ZN(n507) );
  AOI21_X1 U346 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  NAND2_X1 U347 ( .A1(n84), .A2(n85), .ZN(n83) );
  NOR2_X1 U348 ( .A1(n470), .A2(n471), .ZN(n81) );
  OAI211_X1 U350 ( .C1(n436), .C2(n472), .A(n88), .B(n89), .ZN(n82) );
  AND2_X1 U351 ( .A1(n344), .A2(n246), .ZN(n123) );
  OAI21_X1 U353 ( .B1(n14), .B2(n398), .A(n399), .ZN(n344) );
  AND2_X1 U354 ( .A1(n256), .A2(n400), .ZN(n14) );
  AND2_X1 U355 ( .A1(n247), .A2(n244), .ZN(n399) );
  NAND2_X1 U356 ( .A1(n257), .A2(n259), .ZN(n398) );
  NAND2_X1 U357 ( .A1(n121), .A2(n122), .ZN(n77) );
  NAND2_X1 U358 ( .A1(n123), .A2(n124), .ZN(n121) );
  NAND2_X1 U359 ( .A1(n255), .A2(n256), .ZN(n245) );
  NAND2_X1 U360 ( .A1(n257), .A2(n513), .ZN(n255) );
  INV_X1 U361 ( .A(n400), .ZN(n513) );
  INV_X1 U362 ( .A(n259), .ZN(n511) );
  INV_X1 U363 ( .A(n80), .ZN(n469) );
  INV_X1 U364 ( .A(n122), .ZN(n509) );
  OAI211_X1 U365 ( .C1(n285), .C2(n286), .A(n287), .B(n288), .ZN(net497338) );
  NAND4_X1 U366 ( .A1(n304), .A2(net497394), .A3(n305), .A4(n306), .ZN(
        net497232) );
  NAND2_X1 U367 ( .A1(A[11]), .A2(B[11]), .ZN(n338) );
  NAND2_X1 U368 ( .A1(B[12]), .A2(A[12]), .ZN(n325) );
  NOR2_X1 U369 ( .A1(B[17]), .A2(A[17]), .ZN(n1) );
  NOR2_X1 U370 ( .A1(n333), .A2(n53), .ZN(n332) );
  NOR2_X1 U371 ( .A1(A[14]), .A2(B[14]), .ZN(n333) );
  NAND2_X1 U372 ( .A1(B[13]), .A2(A[13]), .ZN(n326) );
  NAND2_X1 U373 ( .A1(A[23]), .A2(B[23]), .ZN(net497316) );
  NAND2_X1 U374 ( .A1(B[29]), .A2(A[29]), .ZN(net497239) );
  NAND2_X1 U375 ( .A1(B[38]), .A2(A[38]), .ZN(net497149) );
  NAND2_X1 U376 ( .A1(B[37]), .A2(A[37]), .ZN(net497154) );
  NAND2_X1 U377 ( .A1(B[62]), .A2(A[62]), .ZN(n85) );
  NAND2_X1 U378 ( .A1(B[53]), .A2(A[53]), .ZN(n143) );
  NAND2_X1 U379 ( .A1(B[57]), .A2(A[57]), .ZN(n112) );
  NAND2_X1 U380 ( .A1(B[61]), .A2(A[61]), .ZN(n88) );
  NAND2_X1 U381 ( .A1(B[54]), .A2(A[54]), .ZN(n144) );
  NAND2_X1 U382 ( .A1(B[58]), .A2(A[58]), .ZN(n113) );
  NAND2_X1 U383 ( .A1(B[49]), .A2(A[49]), .ZN(n178) );
  NAND2_X1 U384 ( .A1(B[56]), .A2(A[56]), .ZN(n111) );
  NAND2_X1 U385 ( .A1(A[15]), .A2(B[15]), .ZN(n318) );
  NAND2_X1 U386 ( .A1(B[60]), .A2(A[60]), .ZN(n89) );
  NAND2_X1 U387 ( .A1(B[45]), .A2(A[45]), .ZN(n206) );
  NAND2_X1 U388 ( .A1(A[8]), .A2(B[8]), .ZN(n63) );
  NAND2_X1 U389 ( .A1(A[18]), .A2(B[18]), .ZN(n306) );
  NAND2_X1 U391 ( .A1(B[14]), .A2(A[14]), .ZN(n346) );
  NAND2_X1 U392 ( .A1(B[10]), .A2(A[10]), .ZN(n377) );
  NAND2_X1 U393 ( .A1(B[36]), .A2(A[36]), .ZN(net497155) );
  NAND2_X1 U394 ( .A1(A[26]), .A2(B[26]), .ZN(n266) );
  NAND2_X1 U395 ( .A1(B[33]), .A2(A[33]), .ZN(net497193) );
  NAND2_X1 U396 ( .A1(B[42]), .A2(A[42]), .ZN(n223) );
  NAND2_X1 U397 ( .A1(B[24]), .A2(A[24]), .ZN(n265) );
  NAND2_X1 U398 ( .A1(B[44]), .A2(A[44]), .ZN(n205) );
  NAND2_X1 U399 ( .A1(B[48]), .A2(A[48]), .ZN(n176) );
  NAND2_X1 U400 ( .A1(B[50]), .A2(A[50]), .ZN(n177) );
  NAND2_X1 U401 ( .A1(B[28]), .A2(A[28]), .ZN(net497238) );
  NAND2_X1 U402 ( .A1(B[6]), .A2(A[6]), .ZN(n66) );
  NAND2_X1 U403 ( .A1(B[52]), .A2(A[52]), .ZN(n142) );
  NAND2_X1 U404 ( .A1(B[46]), .A2(A[46]), .ZN(n207) );
  NAND2_X1 U405 ( .A1(A[19]), .A2(B[19]), .ZN(n305) );
  NAND2_X1 U406 ( .A1(B[41]), .A2(A[41]), .ZN(n227) );
  NAND2_X1 U407 ( .A1(A[27]), .A2(B[27]), .ZN(n274) );
  NAND2_X1 U408 ( .A1(B[32]), .A2(A[32]), .ZN(net497192) );
  NAND2_X1 U409 ( .A1(B[40]), .A2(A[40]), .ZN(n228) );
  NAND2_X1 U410 ( .A1(B[63]), .A2(A[63]), .ZN(n84) );
  INV_X1 U411 ( .A(B[21]), .ZN(n510) );
  NAND2_X1 U412 ( .A1(B[34]), .A2(A[34]), .ZN(net497194) );
  AND2_X1 U413 ( .A1(B[55]), .A2(A[55]), .ZN(n54) );
  AND2_X1 U414 ( .A1(B[59]), .A2(A[59]), .ZN(n55) );
  NAND2_X1 U415 ( .A1(B[47]), .A2(A[47]), .ZN(n191) );
  OR2_X1 U416 ( .A1(B[51]), .A2(A[51]), .ZN(n169) );
  OR2_X1 U417 ( .A1(A[10]), .A2(B[10]), .ZN(n340) );
  OR2_X1 U418 ( .A1(B[63]), .A2(A[63]), .ZN(n80) );
  OR2_X1 U419 ( .A1(B[60]), .A2(A[60]), .ZN(n102) );
  OR2_X1 U420 ( .A1(B[61]), .A2(A[61]), .ZN(n99) );
  OR2_X1 U421 ( .A1(B[62]), .A2(A[62]), .ZN(n95) );
  OR2_X1 U422 ( .A1(A[30]), .A2(B[30]), .ZN(net497243) );
  OR2_X1 U423 ( .A1(B[31]), .A2(A[31]), .ZN(net497244) );
  OR2_X1 U424 ( .A1(B[59]), .A2(A[59]), .ZN(n117) );
  INV_X1 U425 ( .A(B[11]), .ZN(n445) );
  OR2_X1 U426 ( .A1(B[45]), .A2(A[45]), .ZN(n199) );
  OR2_X1 U427 ( .A1(A[8]), .A2(B[8]), .ZN(n62) );
  OR2_X1 U428 ( .A1(B[6]), .A2(A[6]), .ZN(n68) );
  OR2_X1 U429 ( .A1(B[5]), .A2(A[5]), .ZN(n76) );
  OR2_X1 U430 ( .A1(B[2]), .A2(A[2]), .ZN(n259) );
  OR2_X1 U431 ( .A1(B[1]), .A2(A[1]), .ZN(n257) );
  OR2_X1 U432 ( .A1(B[4]), .A2(A[4]), .ZN(n124) );
  OR2_X1 U433 ( .A1(B[3]), .A2(A[3]), .ZN(n246) );
  OR2_X1 U434 ( .A1(B[0]), .A2(A[0]), .ZN(n397) );
  NOR2_X1 U435 ( .A1(n395), .A2(n396), .ZN(n345) );
  NAND2_X1 U436 ( .A1(n68), .A2(n76), .ZN(n395) );
  NAND2_X1 U437 ( .A1(B[4]), .A2(A[4]), .ZN(n122) );
  NAND2_X1 U438 ( .A1(B[1]), .A2(A[1]), .ZN(n256) );
  NAND2_X1 U439 ( .A1(B[2]), .A2(A[2]), .ZN(n244) );
  NAND2_X1 U441 ( .A1(B[0]), .A2(A[0]), .ZN(n400) );
  NAND2_X1 U442 ( .A1(B[5]), .A2(A[5]), .ZN(n75) );
  NAND2_X1 U443 ( .A1(B[3]), .A2(A[3]), .ZN(n247) );
  AND2_X1 U444 ( .A1(A[5]), .A2(B[5]), .ZN(n394) );
  NAND4_X1 U445 ( .A1(net497156), .A2(net497151), .A3(net497153), .A4(
        net497147), .ZN(net497069) );
  OAI21_X1 U446 ( .B1(n11), .B2(net497146), .A(net497147), .ZN(net497068) );
  AOI21_X1 U447 ( .B1(n316), .B2(n9), .A(n312), .ZN(n315) );
  INV_X1 U448 ( .A(net497310), .ZN(n444) );
  NAND2_X1 U449 ( .A1(A[22]), .A2(B[22]), .ZN(n288) );
  OAI21_X1 U450 ( .B1(n443), .B2(net497078), .A(n460), .ZN(net538264) );
  NAND2_X1 U451 ( .A1(n248), .A2(net497194), .ZN(n18) );
  NAND2_X1 U452 ( .A1(net497188), .A2(net497194), .ZN(n249) );
  OAI211_X1 U453 ( .C1(n479), .C2(net497192), .A(net497193), .B(net497194), 
        .ZN(net497190) );
  XNOR2_X1 U454 ( .A(n275), .B(n276), .ZN(SUM[26]) );
  XNOR2_X1 U455 ( .A(n49), .B(n283), .ZN(SUM[24]) );
  AOI21_X1 U456 ( .B1(n497), .B2(n49), .A(n496), .ZN(n275) );
  AND2_X1 U457 ( .A1(n58), .A2(n44), .ZN(n368) );
  NAND2_X1 U458 ( .A1(B[25]), .A2(A[25]), .ZN(n264) );
  NAND2_X1 U459 ( .A1(net497243), .A2(net497240), .ZN(net497267) );
  NAND2_X1 U460 ( .A1(net497250), .A2(net497243), .ZN(net497262) );
  AND2_X1 U461 ( .A1(net497244), .A2(net497243), .ZN(net497233) );
  AND3_X1 U462 ( .A1(net497243), .A2(net497250), .A3(net497249), .ZN(net537151) );
  OAI21_X1 U463 ( .B1(net535589), .B2(n310), .A(n311), .ZN(n309) );
  NAND2_X1 U464 ( .A1(n356), .A2(n326), .ZN(n355) );
  XNOR2_X1 U465 ( .A(n295), .B(net497373), .ZN(SUM[22]) );
  NOR2_X1 U466 ( .A1(A[21]), .A2(B[21]), .ZN(n285) );
  NAND2_X1 U467 ( .A1(B[21]), .A2(A[21]), .ZN(n287) );
  INV_X1 U468 ( .A(A[21]), .ZN(n503) );
  XNOR2_X1 U469 ( .A(n10), .B(n315), .ZN(SUM[18]) );
  NOR2_X1 U470 ( .A1(n485), .A2(n1), .ZN(n320) );
  OAI21_X1 U471 ( .B1(n486), .B2(n1), .A(n314), .ZN(n312) );
  INV_X1 U472 ( .A(n1), .ZN(n484) );
  XNOR2_X1 U473 ( .A(n309), .B(n308), .ZN(SUM[19]) );
  XNOR2_X1 U474 ( .A(n388), .B(n387), .ZN(SUM[10]) );
  OAI21_X1 U475 ( .B1(net537534), .B2(n499), .A(net497239), .ZN(net497268) );
  AND2_X1 U476 ( .A1(net497280), .A2(n41), .ZN(net537534) );
  XNOR2_X1 U477 ( .A(net497267), .B(net497268), .ZN(SUM[30]) );
  AND3_X1 U478 ( .A1(n369), .A2(n368), .A3(n61), .ZN(n39) );
  XNOR2_X1 U479 ( .A(n60), .B(n61), .ZN(SUM[8]) );
  NAND2_X1 U480 ( .A1(n24), .A2(net497153), .ZN(net497167) );
  NAND2_X1 U481 ( .A1(A[35]), .A2(B[35]), .ZN(net497187) );
  OAI21_X1 U482 ( .B1(n136), .B2(n438), .A(n138), .ZN(n134) );
  OAI21_X1 U483 ( .B1(n478), .B2(n438), .A(n142), .ZN(n157) );
  NAND2_X1 U484 ( .A1(n223), .A2(n232), .ZN(n231) );
  NAND2_X1 U485 ( .A1(n318), .A2(n410), .ZN(n347) );
  NAND2_X1 U486 ( .A1(n410), .A2(n351), .ZN(n327) );
  AND2_X1 U487 ( .A1(n410), .A2(n4), .ZN(n2) );
  AND2_X1 U488 ( .A1(n336), .A2(n351), .ZN(n47) );
  NAND2_X1 U489 ( .A1(n282), .A2(n265), .ZN(n281) );
  OAI211_X1 U490 ( .C1(net497311), .C2(n407), .A(n415), .B(n284), .ZN(n49) );
  OAI211_X1 U491 ( .C1(n407), .C2(net497311), .A(net497309), .B(net497312), 
        .ZN(net497310) );
  OAI211_X1 U492 ( .C1(net497311), .C2(n407), .A(net497317), .B(n284), .ZN(
        net497282) );
  AOI21_X1 U493 ( .B1(n342), .B2(n341), .A(n343), .ZN(n329) );
  NAND2_X1 U494 ( .A1(n342), .A2(n372), .ZN(n61) );
  OAI21_X1 U495 ( .B1(n452), .B2(n441), .A(net497154), .ZN(net537813) );
  XNOR2_X1 U496 ( .A(n441), .B(n26), .ZN(SUM[37]) );
  OAI21_X1 U497 ( .B1(n441), .B2(n452), .A(net497154), .ZN(n24) );
  OAI21_X1 U498 ( .B1(n459), .B2(n442), .A(net497155), .ZN(n27) );
  AOI21_X1 U499 ( .B1(n322), .B2(n323), .A(net534733), .ZN(net497441) );
  NOR2_X1 U500 ( .A1(net537101), .A2(n327), .ZN(n322) );
  XNOR2_X1 U501 ( .A(n301), .B(n300), .ZN(SUM[21]) );
  OAI211_X1 U502 ( .C1(n302), .C2(net535589), .A(n286), .B(n296), .ZN(n301) );
  NOR2_X1 U503 ( .A1(n48), .A2(n52), .ZN(n375) );
  NAND2_X1 U504 ( .A1(n364), .A2(n325), .ZN(n363) );
  XNOR2_X1 U505 ( .A(n161), .B(n160), .ZN(SUM[52]) );
  INV_X1 U506 ( .A(n160), .ZN(n438) );
  NAND2_X1 U507 ( .A1(n207), .A2(n210), .ZN(n209) );
  XNOR2_X1 U508 ( .A(net535589), .B(n328), .ZN(SUM[16]) );
  OAI211_X1 U509 ( .C1(n329), .C2(n330), .A(n331), .B(n332), .ZN(n319) );
  AND2_X1 U510 ( .A1(n336), .A2(n4), .ZN(n331) );
  XNOR2_X1 U511 ( .A(net497278), .B(n253), .ZN(SUM[29]) );
  NAND2_X1 U512 ( .A1(n41), .A2(net497280), .ZN(n253) );
  NAND2_X1 U513 ( .A1(n339), .A2(n340), .ZN(n337) );
  NAND2_X1 U514 ( .A1(n389), .A2(n411), .ZN(n388) );
  NAND2_X1 U515 ( .A1(n375), .A2(n339), .ZN(n361) );
  NAND2_X1 U516 ( .A1(n58), .A2(n59), .ZN(n56) );
  AND2_X1 U517 ( .A1(n59), .A2(n63), .ZN(n384) );
  OAI211_X1 U518 ( .C1(n376), .C2(n63), .A(n377), .B(n59), .ZN(n339) );
  INV_X1 U519 ( .A(n27), .ZN(n441) );
  XNOR2_X1 U520 ( .A(net497205), .B(n249), .ZN(SUM[34]) );
  NAND2_X1 U521 ( .A1(B[30]), .A2(A[30]), .ZN(net497240) );
  NAND2_X1 U522 ( .A1(n273), .A2(net497316), .ZN(n272) );
  NAND2_X1 U523 ( .A1(n409), .A2(B[17]), .ZN(n314) );
  XNOR2_X1 U524 ( .A(n158), .B(n157), .ZN(SUM[53]) );
  INV_X1 U525 ( .A(n157), .ZN(n432) );
  NAND2_X1 U526 ( .A1(n162), .A2(n163), .ZN(n160) );
  NAND2_X1 U527 ( .A1(B[51]), .A2(A[51]), .ZN(n174) );
  INV_X1 U528 ( .A(net497190), .ZN(n461) );
  XNOR2_X1 U529 ( .A(n378), .B(n379), .ZN(SUM[11]) );
  NOR2_X1 U531 ( .A1(A[9]), .A2(B[9]), .ZN(n376) );
  NAND2_X1 U532 ( .A1(B[9]), .A2(A[9]), .ZN(n59) );
  NOR2_X1 U533 ( .A1(n443), .A2(net497069), .ZN(net497070) );
  INV_X1 U534 ( .A(net497069), .ZN(n450) );
  NAND2_X1 U535 ( .A1(B[39]), .A2(A[39]), .ZN(net497148) );
  INV_X1 U536 ( .A(net537617), .ZN(n491) );
  AOI211_X1 U537 ( .C1(net497225), .C2(net537617), .A(net537913), .B(n500), 
        .ZN(n31) );
  NAND2_X1 U538 ( .A1(net497282), .A2(net497251), .ZN(n282) );
  AOI21_X1 U539 ( .B1(n481), .B2(net537617), .A(n272), .ZN(net497312) );
  NAND2_X1 U540 ( .A1(net537617), .A2(n481), .ZN(net497317) );
  NAND2_X1 U541 ( .A1(n177), .A2(n181), .ZN(n180) );
  NAND2_X1 U542 ( .A1(n188), .A2(n176), .ZN(n185) );
  NAND2_X1 U543 ( .A1(n17), .A2(net497188), .ZN(n248) );
  OR2_X1 U544 ( .A1(B[47]), .A2(A[47]), .ZN(n201) );
  XNOR2_X1 U545 ( .A(n291), .B(net497359), .ZN(SUM[23]) );
  NAND2_X1 U546 ( .A1(net497348), .A2(n288), .ZN(n295) );
  AND2_X1 U547 ( .A1(net497349), .A2(net497348), .ZN(net497337) );
  AND3_X1 U548 ( .A1(net497349), .A2(net497347), .A3(net497348), .ZN(n290) );
  INV_X1 U549 ( .A(net497348), .ZN(n501) );
  NAND2_X1 U550 ( .A1(n36), .A2(net497348), .ZN(net497366) );
  AND2_X1 U551 ( .A1(n201), .A2(n200), .ZN(n202) );
  XNOR2_X1 U552 ( .A(n57), .B(n56), .ZN(SUM[9]) );
  NAND2_X1 U553 ( .A1(n58), .A2(n57), .ZN(n389) );
  NAND2_X1 U556 ( .A1(n373), .A2(n71), .ZN(n342) );
  OR2_X1 U557 ( .A1(n403), .A2(B[7]), .ZN(n71) );
  OAI21_X1 U558 ( .B1(n403), .B2(B[7]), .A(n124), .ZN(n396) );
  NAND2_X1 U559 ( .A1(A[7]), .A2(B[7]), .ZN(n70) );
  INV_X1 U560 ( .A(n29), .ZN(n442) );
  INV_X1 U561 ( .A(net497143), .ZN(n439) );
  INV_X1 U563 ( .A(n195), .ZN(n457) );
  OAI21_X1 U564 ( .B1(net497062), .B2(n195), .A(n196), .ZN(n194) );
  NAND2_X1 U565 ( .A1(n222), .A2(n221), .ZN(n230) );
  OAI21_X1 U566 ( .B1(n439), .B2(n195), .A(n196), .ZN(n217) );
  OAI21_X1 U567 ( .B1(n219), .B2(n220), .A(n221), .ZN(n196) );
  NAND2_X1 U568 ( .A1(B[43]), .A2(A[43]), .ZN(n222) );
  OAI21_X1 U569 ( .B1(net538090), .B2(n479), .A(net497193), .ZN(net497205) );
  INV_X1 U570 ( .A(n408), .ZN(n443) );
  OAI21_X1 U571 ( .B1(net538090), .B2(n479), .A(net497193), .ZN(n17) );
  NAND2_X1 U572 ( .A1(net497197), .A2(net497195), .ZN(net497212) );
  NAND2_X1 U573 ( .A1(A[31]), .A2(B[31]), .ZN(net497236) );
  OAI21_X1 U575 ( .B1(n443), .B2(net497078), .A(n460), .ZN(n29) );
  INV_X1 U577 ( .A(net497066), .ZN(n460) );
  NAND2_X1 U578 ( .A1(net497188), .A2(net497189), .ZN(net497186) );
  INV_X1 U579 ( .A(n185), .ZN(n431) );
  NAND2_X1 U580 ( .A1(n166), .A2(n167), .ZN(n188) );
  NAND2_X1 U581 ( .A1(n170), .A2(n182), .ZN(n181) );
  XNOR2_X1 U586 ( .A(n233), .B(n234), .ZN(SUM[42]) );
  NAND2_X1 U587 ( .A1(n226), .A2(n233), .ZN(n232) );
  INV_X1 U588 ( .A(n21), .ZN(n440) );
  XNOR2_X1 U591 ( .A(n212), .B(n211), .ZN(SUM[46]) );
  NAND2_X1 U592 ( .A1(n200), .A2(n211), .ZN(n210) );
  NAND2_X1 U593 ( .A1(n217), .A2(n198), .ZN(n216) );
  OAI21_X1 U594 ( .B1(n21), .B2(n458), .A(n227), .ZN(n233) );
  AOI21_X1 U595 ( .B1(n229), .B2(net497143), .A(n455), .ZN(n21) );
  OAI21_X1 U597 ( .B1(n442), .B2(net497069), .A(net497068), .ZN(net497143) );
endmodule


module RCA_NBIT64_13 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_13_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), 
        .SUM({Co, S}) );
endmodule


module RCA_NBIT64_12_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net493900, net493891, net493886, net493885, net493873, net493872,
         net493867, net493866, net493861, net493856, net493845, net493835,
         net493832, net493831, net493830, net493824, net493805, net493791,
         net493788, net493786, net493785, net493779, net537204, net538113,
         net538274, net493850, net493837, net493874, net493871, net493869,
         net493839, net493836, net493887, net493870, net493864, net493858,
         net493841, net493809, net493790, net493865, n2, n3, n8, n9, n10, n11,
         n13, n16, n18, n19, n20, n22, n23, n24, n25, n26, n28, n31, n34, n35,
         n37, n39, n40, n41, n42, n43, n44, n50, n54, n60, n63, n65, n66, n71,
         n74, n75, n76, n78, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90,
         n91, n92, n93, n96, n97, n98, n99, n100, n103, n104, n105, n106, n107,
         n109, n110, n111, n112, n115, n116, n119, n120, n121, n122, n124,
         n125, n126, n128, n129, n130, n131, n132, n133, n134, n136, n137,
         n138, n140, n142, n143, n144, n145, n146, n147, n148, n149, n151,
         n152, n153, n154, n155, n156, n157, n159, n160, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n176,
         n178, n179, n180, n181, n182, n183, n184, n187, n188, n190, n191,
         n192, n193, n194, n195, n196, n197, n200, n201, n202, n204, n205,
         n206, n207, n210, n211, n213, n216, n218, n220, n222, n223, n224,
         n225, n226, n227, n228, n229, n231, n232, n233, n236, n237, n238,
         n239, n240, n241, n242, n243, n245, n247, n248, n249, n251, n252,
         n253, n254, n257, n258, n259, n260, n261, n263, n264, n265, n266,
         n267, n269, n270, n271, n272, n273, n274, n275, n278, n279, n280,
         n281, n282, n283, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n299, n300, n301, n302, n303, n304, n307,
         n308, n309, n310, n314, n315, n316, n317, n318, n320, n323, n324,
         n326, n327, n329, n330, n331, n332, n333, n334, n336, n337, n339,
         n340, n341, n342, n343, n344, n345, n347, n349, n350, n351, n353,
         n354, n356, n357, n358, n359, n360, n361, n362, n363, n364, n367,
         n368, n369, n370, n371, n372, n374, n376, n377, n379, n380, n381,
         n382, n384, n385, n386, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n402, n403, n405, n406, n407, n409, n410,
         n413, n414, n415, n416, n417, n418, n419, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n443, n444, n445, n446, n447, n448, n449,
         n451, n452, n453, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n471, n472, n474, n475, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601;

  OR2_X2 U7 ( .A1(A[33]), .A2(B[33]), .ZN(n273) );
  NAND3_X1 U60 ( .A1(n330), .A2(n357), .A3(n356), .ZN(n329) );
  OR2_X2 U61 ( .A1(B[38]), .A2(A[38]), .ZN(net493871) );
  NOR2_X2 U67 ( .A1(A[9]), .A2(B[9]), .ZN(n86) );
  OR2_X2 U159 ( .A1(B[28]), .A2(A[28]), .ZN(n293) );
  OR2_X2 U160 ( .A1(A[29]), .A2(B[29]), .ZN(n292) );
  OR2_X2 U401 ( .A1(A[22]), .A2(B[22]), .ZN(n303) );
  NAND3_X1 U515 ( .A1(n166), .A2(n167), .A3(n168), .ZN(n165) );
  NAND3_X1 U533 ( .A1(net493779), .A2(n224), .A3(n225), .ZN(n193) );
  NAND3_X1 U556 ( .A1(n3), .A2(n303), .A3(n304), .ZN(n299) );
  NAND3_X1 U563 ( .A1(n334), .A2(n339), .A3(n340), .ZN(n337) );
  NAND3_X1 U567 ( .A1(n332), .A2(n340), .A3(n518), .ZN(n351) );
  NAND3_X1 U568 ( .A1(n303), .A2(n359), .A3(n358), .ZN(n357) );
  NAND3_X1 U575 ( .A1(n390), .A2(n44), .A3(n391), .ZN(n380) );
  NAND3_X1 U584 ( .A1(n446), .A2(n423), .A3(n422), .ZN(n444) );
  NAND3_X1 U585 ( .A1(n452), .A2(n89), .A3(n453), .ZN(n446) );
  OR2_X2 U26 ( .A1(A[10]), .A2(B[10]), .ZN(n426) );
  OR2_X2 U109 ( .A1(B[41]), .A2(A[41]), .ZN(net493836) );
  OR2_X2 U117 ( .A1(B[42]), .A2(A[42]), .ZN(net493837) );
  OR2_X2 U164 ( .A1(B[24]), .A2(A[24]), .ZN(n332) );
  OR2_X2 U165 ( .A1(B[26]), .A2(A[26]), .ZN(n334) );
  OR2_X2 U343 ( .A1(B[46]), .A2(A[46]), .ZN(n236) );
  OR2_X2 U364 ( .A1(B[34]), .A2(A[34]), .ZN(n265) );
  CLKBUF_X1 U2 ( .A(n78), .Z(n478) );
  INV_X1 U3 ( .A(n574), .ZN(n479) );
  INV_X1 U4 ( .A(n492), .ZN(n389) );
  OR2_X1 U5 ( .A1(B[12]), .A2(A[12]), .ZN(n414) );
  OR2_X1 U6 ( .A1(A[17]), .A2(B[17]), .ZN(n385) );
  OR2_X1 U8 ( .A1(A[27]), .A2(B[27]), .ZN(n490) );
  AND2_X1 U9 ( .A1(n394), .A2(n475), .ZN(SUM[0]) );
  OR2_X1 U10 ( .A1(B[32]), .A2(A[32]), .ZN(n272) );
  NOR2_X1 U11 ( .A1(A[30]), .A2(B[30]), .ZN(n13) );
  OR2_X1 U12 ( .A1(B[36]), .A2(A[36]), .ZN(net493874) );
  OR2_X1 U13 ( .A1(B[44]), .A2(A[44]), .ZN(n238) );
  OR2_X1 U14 ( .A1(B[40]), .A2(A[40]), .ZN(net493841) );
  OR2_X1 U15 ( .A1(B[43]), .A2(A[43]), .ZN(net493831) );
  OR2_X1 U16 ( .A1(B[37]), .A2(A[37]), .ZN(net493869) );
  OR2_X1 U17 ( .A1(A[35]), .A2(B[35]), .ZN(n266) );
  OR2_X1 U18 ( .A1(B[45]), .A2(A[45]), .ZN(n239) );
  OR2_X1 U19 ( .A1(B[49]), .A2(A[49]), .ZN(n216) );
  OR2_X1 U20 ( .A1(B[48]), .A2(A[48]), .ZN(n200) );
  OR2_X1 U21 ( .A1(B[50]), .A2(A[50]), .ZN(n196) );
  AND2_X1 U22 ( .A1(n513), .A2(n514), .ZN(n187) );
  OR2_X1 U23 ( .A1(B[53]), .A2(A[53]), .ZN(n172) );
  OR2_X1 U24 ( .A1(B[54]), .A2(A[54]), .ZN(n169) );
  OR2_X1 U25 ( .A1(B[55]), .A2(A[55]), .ZN(n170) );
  OR2_X1 U27 ( .A1(B[52]), .A2(A[52]), .ZN(n171) );
  OR2_X1 U28 ( .A1(B[56]), .A2(A[56]), .ZN(n147) );
  OR2_X1 U29 ( .A1(B[57]), .A2(A[57]), .ZN(n148) );
  OR2_X1 U30 ( .A1(B[58]), .A2(A[58]), .ZN(n145) );
  CLKBUF_X1 U31 ( .A(n314), .Z(n480) );
  NOR2_X1 U32 ( .A1(B[47]), .A2(A[47]), .ZN(n481) );
  AND2_X1 U33 ( .A1(A[18]), .A2(B[18]), .ZN(n482) );
  CLKBUF_X1 U34 ( .A(A[18]), .Z(n483) );
  CLKBUF_X1 U35 ( .A(n337), .Z(n484) );
  OR2_X2 U36 ( .A1(B[25]), .A2(A[25]), .ZN(n333) );
  CLKBUF_X1 U37 ( .A(net493788), .Z(n485) );
  XNOR2_X1 U38 ( .A(n18), .B(n438), .ZN(SUM[15]) );
  INV_X1 U39 ( .A(n490), .ZN(n486) );
  NAND4_X1 U40 ( .A1(n490), .A2(n333), .A3(n334), .A4(n332), .ZN(n487) );
  OAI21_X1 U41 ( .B1(n497), .B2(net493809), .A(net493790), .ZN(n488) );
  BUF_X1 U42 ( .A(n341), .Z(n489) );
  XNOR2_X1 U43 ( .A(n499), .B(n491), .ZN(SUM[49]) );
  NAND2_X1 U44 ( .A1(n222), .A2(n205), .ZN(n491) );
  AND2_X2 U45 ( .A1(B[16]), .A2(A[16]), .ZN(n492) );
  NAND2_X1 U46 ( .A1(n386), .A2(n482), .ZN(n379) );
  AND2_X1 U47 ( .A1(n249), .A2(n231), .ZN(n493) );
  NAND2_X1 U48 ( .A1(n364), .A2(n367), .ZN(n494) );
  OR2_X2 U49 ( .A1(B[51]), .A2(A[51]), .ZN(n197) );
  OR2_X1 U50 ( .A1(A[19]), .A2(B[19]), .ZN(n44) );
  XNOR2_X1 U51 ( .A(n495), .B(n497), .ZN(SUM[36]) );
  AND2_X1 U52 ( .A1(net493874), .A2(net493873), .ZN(n495) );
  XNOR2_X1 U53 ( .A(n66), .B(n496), .ZN(SUM[35]) );
  NAND2_X1 U54 ( .A1(n264), .A2(n266), .ZN(n496) );
  CLKBUF_X1 U55 ( .A(n16), .Z(n497) );
  XOR2_X1 U56 ( .A(n498), .B(n374), .Z(SUM[21]) );
  NAND2_X1 U57 ( .A1(n494), .A2(n361), .ZN(n498) );
  NAND2_X1 U58 ( .A1(n216), .A2(n206), .ZN(n499) );
  XOR2_X1 U59 ( .A(n500), .B(n532), .Z(SUM[33]) );
  AND2_X1 U62 ( .A1(n273), .A2(n270), .ZN(n500) );
  XOR2_X1 U63 ( .A(n20), .B(n501), .Z(SUM[25]) );
  NAND2_X1 U64 ( .A1(n342), .A2(n353), .ZN(n501) );
  XNOR2_X1 U65 ( .A(n502), .B(n354), .ZN(SUM[24]) );
  NAND2_X1 U66 ( .A1(n332), .A2(n342), .ZN(n502) );
  XOR2_X1 U68 ( .A(n503), .B(net538113), .Z(SUM[32]) );
  AND2_X1 U69 ( .A1(n272), .A2(n269), .ZN(n503) );
  XOR2_X1 U70 ( .A(n504), .B(n184), .Z(SUM[54]) );
  AND2_X1 U71 ( .A1(n169), .A2(n179), .ZN(n504) );
  XOR2_X1 U72 ( .A(n520), .B(n505), .Z(SUM[30]) );
  AND2_X1 U73 ( .A1(n581), .A2(n287), .ZN(n505) );
  AOI21_X1 U74 ( .B1(n570), .B2(net538113), .A(net493788), .ZN(n16) );
  INV_X1 U75 ( .A(net493805), .ZN(n570) );
  XNOR2_X1 U76 ( .A(n326), .B(n327), .ZN(SUM[28]) );
  NOR2_X1 U77 ( .A1(n577), .A2(n578), .ZN(n327) );
  NOR2_X1 U78 ( .A1(n23), .A2(n519), .ZN(n326) );
  INV_X1 U79 ( .A(n323), .ZN(n519) );
  XNOR2_X1 U80 ( .A(n523), .B(n261), .ZN(SUM[37]) );
  NOR2_X1 U81 ( .A1(n567), .A2(n566), .ZN(n261) );
  INV_X1 U82 ( .A(n132), .ZN(n528) );
  NAND2_X1 U83 ( .A1(n357), .A2(n356), .ZN(n331) );
  INV_X1 U84 ( .A(n299), .ZN(n540) );
  OR2_X1 U85 ( .A1(n296), .A2(n65), .ZN(n323) );
  NAND2_X1 U86 ( .A1(n336), .A2(n329), .ZN(n65) );
  INV_X1 U87 ( .A(n43), .ZN(n535) );
  OAI21_X1 U88 ( .B1(n80), .B2(n429), .A(n464), .ZN(n89) );
  AOI21_X1 U89 ( .B1(n106), .B2(n107), .A(n550), .ZN(SUM[64]) );
  XNOR2_X1 U90 ( .A(n8), .B(n405), .ZN(SUM[17]) );
  NAND2_X1 U91 ( .A1(n402), .A2(n385), .ZN(n405) );
  NAND2_X1 U92 ( .A1(n406), .A2(n389), .ZN(n8) );
  NAND2_X1 U93 ( .A1(n389), .A2(n392), .ZN(n407) );
  AOI21_X1 U94 ( .B1(n137), .B2(n138), .A(n548), .ZN(n136) );
  NAND4_X1 U95 ( .A1(n147), .A2(n148), .A3(n145), .A4(n146), .ZN(n134) );
  OAI211_X1 U96 ( .C1(n549), .C2(n142), .A(n143), .B(n144), .ZN(n138) );
  NAND2_X1 U97 ( .A1(n432), .A2(n437), .ZN(n440) );
  NAND2_X1 U98 ( .A1(n421), .A2(n413), .ZN(n438) );
  NAND2_X1 U99 ( .A1(n334), .A2(n343), .ZN(n349) );
  NAND2_X1 U100 ( .A1(n423), .A2(n451), .ZN(n458) );
  NAND2_X1 U101 ( .A1(n414), .A2(n435), .ZN(n445) );
  NAND2_X1 U102 ( .A1(net493837), .A2(n41), .ZN(net493850) );
  NAND2_X1 U103 ( .A1(n44), .A2(n382), .ZN(n395) );
  NAND2_X1 U104 ( .A1(n205), .A2(n200), .ZN(n223) );
  NAND2_X1 U105 ( .A1(net493841), .A2(n37), .ZN(net493861) );
  XOR2_X1 U106 ( .A(n506), .B(n480), .Z(SUM[29]) );
  AND2_X1 U107 ( .A1(n286), .A2(n292), .ZN(n506) );
  XOR2_X1 U108 ( .A(n507), .B(n213), .Z(SUM[50]) );
  AND2_X1 U110 ( .A1(n196), .A2(n207), .ZN(n507) );
  XOR2_X1 U111 ( .A(n508), .B(net493824), .Z(SUM[44]) );
  AND2_X1 U112 ( .A1(n238), .A2(n231), .ZN(n508) );
  NAND2_X1 U113 ( .A1(n147), .A2(n142), .ZN(n163) );
  NAND2_X1 U114 ( .A1(n148), .A2(n143), .ZN(n160) );
  NAND2_X1 U115 ( .A1(n265), .A2(n271), .ZN(n275) );
  NAND2_X1 U116 ( .A1(n426), .A2(n449), .ZN(n462) );
  NAND2_X1 U118 ( .A1(n26), .A2(n363), .ZN(n369) );
  NAND2_X1 U119 ( .A1(n370), .A2(n303), .ZN(n26) );
  INV_X1 U120 ( .A(n147), .ZN(n554) );
  NOR2_X1 U121 ( .A1(n538), .A2(n539), .ZN(n374) );
  INV_X1 U122 ( .A(n360), .ZN(n538) );
  INV_X1 U123 ( .A(n269), .ZN(n568) );
  INV_X1 U124 ( .A(n37), .ZN(n558) );
  INV_X1 U125 ( .A(n286), .ZN(n582) );
  OAI211_X1 U126 ( .C1(n545), .C2(n205), .A(n206), .B(n207), .ZN(n202) );
  INV_X1 U127 ( .A(n204), .ZN(n543) );
  OAI21_X1 U128 ( .B1(n529), .B2(n549), .A(n143), .ZN(n156) );
  OAI21_X1 U129 ( .B1(n528), .B2(n553), .A(n116), .ZN(n129) );
  OAI21_X1 U130 ( .B1(n527), .B2(n552), .A(n115), .ZN(n125) );
  INV_X1 U131 ( .A(n129), .ZN(n527) );
  NAND4_X1 U132 ( .A1(n279), .A2(n278), .A3(n280), .A4(n281), .ZN(net538113)
         );
  NAND2_X1 U133 ( .A1(net493836), .A2(net493839), .ZN(net493856) );
  OAI21_X1 U134 ( .B1(n559), .B2(n522), .A(n37), .ZN(net538274) );
  INV_X1 U135 ( .A(net493841), .ZN(n559) );
  NOR2_X1 U136 ( .A1(n481), .A2(n82), .ZN(n242) );
  INV_X1 U137 ( .A(n233), .ZN(n563) );
  AND3_X1 U138 ( .A1(net493869), .A2(net493870), .A3(net493871), .ZN(n9) );
  NAND2_X1 U139 ( .A1(net493872), .A2(net493873), .ZN(net493870) );
  NAND2_X1 U140 ( .A1(net493871), .A2(net493867), .ZN(net493891) );
  INV_X1 U141 ( .A(net493874), .ZN(n555) );
  AND2_X1 U142 ( .A1(net493839), .A2(n37), .ZN(n10) );
  XNOR2_X1 U143 ( .A(n133), .B(n132), .ZN(SUM[60]) );
  NAND2_X1 U144 ( .A1(n131), .A2(n116), .ZN(n133) );
  OAI21_X1 U145 ( .B1(n525), .B2(n547), .A(n180), .ZN(n184) );
  INV_X1 U146 ( .A(n187), .ZN(n525) );
  AOI21_X1 U147 ( .B1(n573), .B2(n484), .A(n575), .ZN(n23) );
  OAI21_X1 U148 ( .B1(n493), .B2(n564), .A(n232), .ZN(n243) );
  XNOR2_X1 U149 ( .A(n377), .B(n60), .ZN(SUM[20]) );
  NAND2_X1 U150 ( .A1(n367), .A2(n361), .ZN(n377) );
  XNOR2_X1 U151 ( .A(n190), .B(n168), .ZN(SUM[52]) );
  NAND2_X1 U152 ( .A1(n171), .A2(n178), .ZN(n190) );
  XNOR2_X1 U153 ( .A(n370), .B(n371), .ZN(SUM[22]) );
  NAND2_X1 U154 ( .A1(n363), .A2(n303), .ZN(n371) );
  XNOR2_X1 U155 ( .A(n248), .B(n247), .ZN(SUM[45]) );
  NAND2_X1 U156 ( .A1(n239), .A2(n232), .ZN(n248) );
  XNOR2_X1 U157 ( .A(n157), .B(n156), .ZN(SUM[58]) );
  NAND2_X1 U158 ( .A1(n145), .A2(n144), .ZN(n157) );
  XNOR2_X1 U161 ( .A(n130), .B(n129), .ZN(SUM[61]) );
  NAND2_X1 U162 ( .A1(n128), .A2(n115), .ZN(n130) );
  XNOR2_X1 U163 ( .A(n126), .B(n125), .ZN(SUM[62]) );
  NAND2_X1 U166 ( .A1(n124), .A2(n120), .ZN(n126) );
  XNOR2_X1 U167 ( .A(n243), .B(n245), .ZN(SUM[46]) );
  NAND2_X1 U168 ( .A1(n236), .A2(n233), .ZN(n245) );
  XNOR2_X1 U169 ( .A(n517), .B(n399), .ZN(SUM[18]) );
  NOR2_X1 U170 ( .A1(n403), .A2(n537), .ZN(n399) );
  INV_X1 U171 ( .A(n397), .ZN(n537) );
  AND2_X1 U172 ( .A1(n489), .A2(n340), .ZN(n20) );
  NAND2_X1 U173 ( .A1(n354), .A2(n332), .ZN(n353) );
  NAND2_X1 U174 ( .A1(n561), .A2(n226), .ZN(n225) );
  OAI21_X1 U175 ( .B1(n569), .B2(n263), .A(n264), .ZN(net493788) );
  OAI211_X1 U176 ( .C1(n571), .C2(n269), .A(n270), .B(n271), .ZN(n267) );
  AOI21_X1 U177 ( .B1(n573), .B2(n337), .A(n486), .ZN(n289) );
  NAND4_X1 U178 ( .A1(n3), .A2(n303), .A3(n304), .A4(n60), .ZN(n330) );
  OAI211_X1 U179 ( .C1(n417), .C2(n418), .A(n414), .B(n419), .ZN(n410) );
  AOI21_X1 U180 ( .B1(n464), .B2(n424), .A(n416), .ZN(n417) );
  NAND2_X1 U181 ( .A1(n2), .A2(n423), .ZN(n418) );
  XNOR2_X1 U182 ( .A(n121), .B(n122), .ZN(SUM[63]) );
  NAND2_X1 U183 ( .A1(n119), .A2(n109), .ZN(n121) );
  OAI21_X1 U184 ( .B1(n526), .B2(n551), .A(n120), .ZN(n122) );
  INV_X1 U185 ( .A(n125), .ZN(n526) );
  OAI21_X1 U186 ( .B1(n512), .B2(n545), .A(n206), .ZN(n213) );
  OAI21_X1 U187 ( .B1(n76), .B2(n534), .A(n436), .ZN(n439) );
  NAND4_X1 U188 ( .A1(n44), .A2(n385), .A3(n392), .A4(n390), .ZN(n307) );
  XNOR2_X1 U189 ( .A(n188), .B(n187), .ZN(SUM[53]) );
  NAND2_X1 U190 ( .A1(n172), .A2(n180), .ZN(n188) );
  XNOR2_X1 U191 ( .A(net493886), .B(net493885), .ZN(SUM[39]) );
  NAND2_X1 U192 ( .A1(net493887), .A2(net493867), .ZN(net493886) );
  NAND2_X1 U193 ( .A1(n524), .A2(net493871), .ZN(net493887) );
  XNOR2_X1 U194 ( .A(n309), .B(n310), .ZN(SUM[31]) );
  NOR2_X1 U195 ( .A1(n478), .A2(n580), .ZN(n310) );
  NAND2_X1 U196 ( .A1(n24), .A2(n25), .ZN(n309) );
  INV_X1 U197 ( .A(n281), .ZN(n580) );
  NOR2_X1 U198 ( .A1(n585), .A2(n584), .ZN(n453) );
  OAI211_X1 U199 ( .C1(n583), .C2(n285), .A(n286), .B(n287), .ZN(n283) );
  NOR2_X1 U200 ( .A1(n78), .A2(n13), .ZN(n282) );
  INV_X1 U201 ( .A(n292), .ZN(n583) );
  OAI211_X1 U202 ( .C1(n564), .C2(n231), .A(n232), .B(n233), .ZN(n229) );
  NAND4_X1 U203 ( .A1(n240), .A2(n239), .A3(n236), .A4(n238), .ZN(net493791)
         );
  NAND2_X1 U204 ( .A1(n595), .A2(n572), .ZN(n336) );
  NAND4_X1 U205 ( .A1(n302), .A2(n300), .A3(n301), .A4(n581), .ZN(n278) );
  NOR2_X1 U206 ( .A1(n78), .A2(n299), .ZN(n302) );
  INV_X1 U207 ( .A(n490), .ZN(n575) );
  INV_X1 U208 ( .A(n216), .ZN(n545) );
  NOR2_X1 U209 ( .A1(n545), .A2(n541), .ZN(n195) );
  INV_X1 U210 ( .A(n200), .ZN(n541) );
  AOI21_X1 U211 ( .B1(n173), .B2(n174), .A(n546), .ZN(n164) );
  OAI211_X1 U212 ( .C1(n547), .C2(n178), .A(n179), .B(n180), .ZN(n174) );
  AOI21_X1 U213 ( .B1(n294), .B2(n295), .A(n296), .ZN(n288) );
  NOR2_X1 U214 ( .A1(n291), .A2(n78), .ZN(n290) );
  NAND2_X1 U215 ( .A1(n540), .A2(n535), .ZN(n295) );
  NAND2_X1 U216 ( .A1(n595), .A2(n572), .ZN(n304) );
  NAND2_X1 U217 ( .A1(n176), .A2(n170), .ZN(n181) );
  NOR2_X1 U218 ( .A1(n481), .A2(n562), .ZN(n228) );
  INV_X1 U219 ( .A(n236), .ZN(n562) );
  OR2_X1 U220 ( .A1(n579), .A2(n342), .ZN(n22) );
  INV_X1 U221 ( .A(n13), .ZN(n581) );
  AND2_X1 U222 ( .A1(n463), .A2(n91), .ZN(n83) );
  NAND2_X1 U223 ( .A1(n89), .A2(n90), .ZN(n463) );
  NAND2_X1 U224 ( .A1(n287), .A2(n13), .ZN(n25) );
  INV_X1 U225 ( .A(n131), .ZN(n553) );
  INV_X1 U226 ( .A(n128), .ZN(n552) );
  INV_X1 U227 ( .A(n124), .ZN(n551) );
  INV_X1 U228 ( .A(n239), .ZN(n564) );
  INV_X1 U229 ( .A(n148), .ZN(n549) );
  INV_X1 U230 ( .A(n172), .ZN(n547) );
  NAND2_X1 U231 ( .A1(n421), .A2(n54), .ZN(n409) );
  INV_X1 U232 ( .A(net493872), .ZN(n567) );
  INV_X1 U233 ( .A(n293), .ZN(n578) );
  XNOR2_X1 U234 ( .A(n153), .B(n154), .ZN(SUM[59]) );
  NAND2_X1 U235 ( .A1(n140), .A2(n146), .ZN(n153) );
  NAND2_X1 U236 ( .A1(n155), .A2(n144), .ZN(n154) );
  NAND2_X1 U237 ( .A1(n145), .A2(n156), .ZN(n155) );
  INV_X1 U238 ( .A(net493869), .ZN(n566) );
  INV_X1 U239 ( .A(n285), .ZN(n577) );
  INV_X1 U240 ( .A(n273), .ZN(n571) );
  AND2_X1 U241 ( .A1(n426), .A2(n451), .ZN(n447) );
  NAND2_X1 U242 ( .A1(n341), .A2(n342), .ZN(n339) );
  NAND2_X1 U243 ( .A1(n360), .A2(n361), .ZN(n359) );
  OAI21_X1 U244 ( .B1(n74), .B2(n536), .A(n402), .ZN(n398) );
  INV_X1 U245 ( .A(n385), .ZN(n536) );
  AND2_X1 U246 ( .A1(n406), .A2(n389), .ZN(n74) );
  INV_X1 U247 ( .A(n176), .ZN(n546) );
  NAND2_X1 U248 ( .A1(net493836), .A2(net493837), .ZN(net493835) );
  INV_X1 U249 ( .A(net493836), .ZN(n565) );
  AND2_X1 U250 ( .A1(n146), .A2(n145), .ZN(n137) );
  OAI21_X1 U251 ( .B1(n372), .B2(n539), .A(n360), .ZN(n370) );
  AND2_X1 U252 ( .A1(n376), .A2(n361), .ZN(n372) );
  AND2_X1 U253 ( .A1(n170), .A2(n169), .ZN(n173) );
  INV_X1 U254 ( .A(n196), .ZN(n544) );
  INV_X1 U255 ( .A(n140), .ZN(n548) );
  INV_X1 U256 ( .A(n343), .ZN(n576) );
  AND2_X1 U257 ( .A1(n169), .A2(n170), .ZN(n167) );
  AND2_X1 U258 ( .A1(n171), .A2(n172), .ZN(n166) );
  XNOR2_X1 U259 ( .A(n83), .B(n84), .ZN(SUM[9]) );
  INV_X1 U260 ( .A(n87), .ZN(n586) );
  XNOR2_X1 U261 ( .A(n393), .B(n601), .ZN(SUM[1]) );
  NAND2_X1 U262 ( .A1(n318), .A2(n317), .ZN(n393) );
  XNOR2_X1 U263 ( .A(n149), .B(n104), .ZN(SUM[5]) );
  NAND2_X1 U264 ( .A1(n152), .A2(n103), .ZN(n149) );
  XNOR2_X1 U265 ( .A(n100), .B(n97), .ZN(SUM[6]) );
  NAND2_X1 U266 ( .A1(n105), .A2(n96), .ZN(n100) );
  XNOR2_X1 U267 ( .A(n88), .B(n89), .ZN(SUM[8]) );
  NAND2_X1 U268 ( .A1(n90), .A2(n91), .ZN(n88) );
  XNOR2_X1 U269 ( .A(n80), .B(n218), .ZN(SUM[4]) );
  NOR2_X1 U270 ( .A1(n594), .A2(n593), .ZN(n218) );
  INV_X1 U271 ( .A(n151), .ZN(n594) );
  INV_X1 U272 ( .A(n220), .ZN(n593) );
  XNOR2_X1 U273 ( .A(n92), .B(n93), .ZN(SUM[7]) );
  OAI21_X1 U274 ( .B1(n590), .B2(n589), .A(n96), .ZN(n93) );
  NAND2_X1 U275 ( .A1(n98), .A2(n99), .ZN(n92) );
  INV_X1 U276 ( .A(n97), .ZN(n590) );
  XNOR2_X1 U277 ( .A(n315), .B(n258), .ZN(SUM[2]) );
  NAND2_X1 U278 ( .A1(n320), .A2(n257), .ZN(n315) );
  XNOR2_X1 U279 ( .A(n253), .B(n254), .ZN(SUM[3]) );
  OAI21_X1 U280 ( .B1(n599), .B2(n598), .A(n257), .ZN(n254) );
  NAND2_X1 U281 ( .A1(n259), .A2(n260), .ZN(n253) );
  INV_X1 U282 ( .A(n258), .ZN(n599) );
  OAI21_X1 U283 ( .B1(n593), .B2(n80), .A(n151), .ZN(n104) );
  OAI21_X1 U284 ( .B1(n592), .B2(n591), .A(n103), .ZN(n97) );
  INV_X1 U285 ( .A(n104), .ZN(n592) );
  AND2_X1 U286 ( .A1(n99), .A2(n465), .ZN(n464) );
  OAI21_X1 U287 ( .B1(n466), .B2(n467), .A(n468), .ZN(n465) );
  NAND4_X1 U288 ( .A1(n220), .A2(n152), .A3(n105), .A4(n98), .ZN(n429) );
  OAI21_X1 U289 ( .B1(n600), .B2(n471), .A(n472), .ZN(n428) );
  INV_X1 U290 ( .A(n474), .ZN(n600) );
  NAND2_X1 U291 ( .A1(n257), .A2(n317), .ZN(n471) );
  NOR2_X1 U292 ( .A1(n597), .A2(n598), .ZN(n472) );
  OAI21_X1 U293 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  NAND2_X1 U294 ( .A1(n115), .A2(n116), .ZN(n111) );
  NOR2_X1 U295 ( .A1(n528), .A2(n553), .ZN(n110) );
  NOR2_X1 U296 ( .A1(n551), .A2(n552), .ZN(n112) );
  AND2_X1 U297 ( .A1(n260), .A2(n428), .ZN(n80) );
  INV_X1 U298 ( .A(n90), .ZN(n587) );
  NOR2_X1 U299 ( .A1(n588), .A2(n589), .ZN(n468) );
  INV_X1 U300 ( .A(n98), .ZN(n588) );
  NAND2_X1 U301 ( .A1(n316), .A2(n317), .ZN(n258) );
  NAND2_X1 U302 ( .A1(n318), .A2(n601), .ZN(n316) );
  NOR2_X1 U303 ( .A1(n591), .A2(n151), .ZN(n466) );
  INV_X1 U304 ( .A(n394), .ZN(n601) );
  INV_X1 U305 ( .A(n105), .ZN(n589) );
  INV_X1 U306 ( .A(n152), .ZN(n591) );
  INV_X1 U307 ( .A(n320), .ZN(n598) );
  NAND2_X1 U308 ( .A1(n96), .A2(n103), .ZN(n467) );
  OR2_X1 U309 ( .A1(n429), .A2(n81), .ZN(n424) );
  AND2_X1 U310 ( .A1(n428), .A2(n260), .ZN(n81) );
  INV_X1 U311 ( .A(n426), .ZN(n585) );
  AND2_X1 U312 ( .A1(n119), .A2(n120), .ZN(n106) );
  INV_X1 U313 ( .A(n427), .ZN(n584) );
  INV_X1 U314 ( .A(n259), .ZN(n597) );
  INV_X1 U315 ( .A(n109), .ZN(n550) );
  NOR2_X1 U316 ( .A1(n11), .A2(n575), .ZN(n345) );
  XOR2_X1 U317 ( .A(n509), .B(n441), .Z(SUM[13]) );
  AND2_X1 U318 ( .A1(n415), .A2(n436), .ZN(n509) );
  NAND2_X1 U319 ( .A1(A[30]), .A2(B[30]), .ZN(n287) );
  NAND2_X1 U320 ( .A1(B[40]), .A2(A[40]), .ZN(n37) );
  NAND2_X1 U321 ( .A1(B[24]), .A2(A[24]), .ZN(n342) );
  OR2_X1 U322 ( .A1(B[18]), .A2(A[18]), .ZN(n390) );
  NAND2_X1 U323 ( .A1(B[20]), .A2(A[20]), .ZN(n361) );
  NAND2_X1 U324 ( .A1(B[53]), .A2(A[53]), .ZN(n180) );
  NAND2_X1 U325 ( .A1(A[31]), .A2(B[31]), .ZN(n281) );
  NAND2_X1 U326 ( .A1(B[58]), .A2(A[58]), .ZN(n144) );
  NAND2_X1 U327 ( .A1(B[60]), .A2(A[60]), .ZN(n116) );
  NAND2_X1 U328 ( .A1(B[32]), .A2(A[32]), .ZN(n269) );
  NAND2_X1 U329 ( .A1(B[46]), .A2(A[46]), .ZN(n233) );
  NAND2_X1 U330 ( .A1(B[57]), .A2(A[57]), .ZN(n143) );
  NAND2_X1 U331 ( .A1(B[52]), .A2(A[52]), .ZN(n178) );
  NAND2_X1 U332 ( .A1(B[49]), .A2(A[49]), .ZN(n206) );
  NAND2_X1 U333 ( .A1(B[45]), .A2(A[45]), .ZN(n232) );
  NAND2_X1 U334 ( .A1(B[26]), .A2(A[26]), .ZN(n343) );
  NAND2_X1 U335 ( .A1(B[12]), .A2(A[12]), .ZN(n435) );
  NAND2_X1 U336 ( .A1(B[61]), .A2(A[61]), .ZN(n115) );
  NAND2_X1 U337 ( .A1(B[29]), .A2(A[29]), .ZN(n286) );
  NAND2_X1 U338 ( .A1(B[21]), .A2(A[21]), .ZN(n360) );
  NAND2_X1 U339 ( .A1(B[41]), .A2(A[41]), .ZN(net493839) );
  NAND2_X1 U340 ( .A1(B[44]), .A2(A[44]), .ZN(n231) );
  NAND2_X1 U341 ( .A1(B[56]), .A2(A[56]), .ZN(n142) );
  NAND2_X1 U342 ( .A1(B[38]), .A2(A[38]), .ZN(net493867) );
  NAND2_X1 U344 ( .A1(B[36]), .A2(A[36]), .ZN(net493873) );
  NAND2_X1 U345 ( .A1(A[22]), .A2(B[22]), .ZN(n363) );
  NAND2_X1 U346 ( .A1(B[54]), .A2(A[54]), .ZN(n179) );
  NAND2_X1 U347 ( .A1(B[62]), .A2(A[62]), .ZN(n120) );
  NAND2_X1 U348 ( .A1(B[34]), .A2(A[34]), .ZN(n271) );
  NAND2_X1 U349 ( .A1(B[50]), .A2(A[50]), .ZN(n207) );
  NAND2_X1 U350 ( .A1(B[37]), .A2(A[37]), .ZN(net493872) );
  NAND2_X1 U351 ( .A1(B[9]), .A2(A[9]), .ZN(n87) );
  OAI21_X1 U352 ( .B1(n574), .B2(n596), .A(n343), .ZN(n31) );
  INV_X1 U353 ( .A(B[27]), .ZN(n596) );
  NAND2_X1 U354 ( .A1(B[42]), .A2(A[42]), .ZN(n41) );
  OR2_X1 U355 ( .A1(B[59]), .A2(A[59]), .ZN(n146) );
  NAND2_X1 U356 ( .A1(B[15]), .A2(A[15]), .ZN(n413) );
  OR2_X1 U357 ( .A1(B[16]), .A2(A[16]), .ZN(n392) );
  NAND2_X1 U358 ( .A1(B[17]), .A2(A[17]), .ZN(n402) );
  NAND2_X1 U359 ( .A1(B[28]), .A2(A[28]), .ZN(n285) );
  NAND2_X1 U360 ( .A1(B[59]), .A2(A[59]), .ZN(n140) );
  AND2_X1 U361 ( .A1(A[17]), .A2(B[17]), .ZN(n391) );
  NAND2_X1 U362 ( .A1(A[35]), .A2(B[35]), .ZN(n264) );
  OR2_X1 U363 ( .A1(A[15]), .A2(B[15]), .ZN(n421) );
  NAND2_X1 U365 ( .A1(B[51]), .A2(A[51]), .ZN(n204) );
  INV_X1 U366 ( .A(B[23]), .ZN(n595) );
  NAND2_X1 U367 ( .A1(B[63]), .A2(A[63]), .ZN(n119) );
  OR2_X1 U368 ( .A1(B[47]), .A2(A[47]), .ZN(n240) );
  OR2_X1 U369 ( .A1(B[63]), .A2(A[63]), .ZN(n109) );
  OR2_X1 U370 ( .A1(B[60]), .A2(A[60]), .ZN(n131) );
  OR2_X1 U371 ( .A1(B[61]), .A2(A[61]), .ZN(n128) );
  OR2_X1 U372 ( .A1(B[62]), .A2(A[62]), .ZN(n124) );
  NAND2_X1 U373 ( .A1(n510), .A2(n511), .ZN(n291) );
  OR2_X1 U374 ( .A1(B[30]), .A2(A[30]), .ZN(n510) );
  AND2_X1 U375 ( .A1(n292), .A2(n293), .ZN(n511) );
  OR2_X1 U376 ( .A1(B[20]), .A2(A[20]), .ZN(n367) );
  OR2_X1 U377 ( .A1(A[39]), .A2(B[39]), .ZN(net493865) );
  OR2_X1 U378 ( .A1(A[21]), .A2(B[21]), .ZN(n358) );
  OR2_X1 U379 ( .A1(B[13]), .A2(A[13]), .ZN(n415) );
  INV_X1 U380 ( .A(n433), .ZN(n533) );
  OAI211_X1 U381 ( .C1(n434), .C2(n435), .A(n436), .B(n437), .ZN(n433) );
  NOR2_X1 U382 ( .A1(A[31]), .A2(B[31]), .ZN(n78) );
  OR2_X1 U383 ( .A1(B[8]), .A2(A[8]), .ZN(n90) );
  OR2_X1 U384 ( .A1(B[7]), .A2(A[7]), .ZN(n98) );
  OR2_X1 U385 ( .A1(B[6]), .A2(A[6]), .ZN(n105) );
  OR2_X1 U386 ( .A1(B[5]), .A2(A[5]), .ZN(n152) );
  OR2_X1 U387 ( .A1(B[2]), .A2(A[2]), .ZN(n320) );
  OR2_X1 U388 ( .A1(B[3]), .A2(A[3]), .ZN(n259) );
  OR2_X1 U389 ( .A1(B[1]), .A2(A[1]), .ZN(n318) );
  OR2_X1 U390 ( .A1(B[4]), .A2(A[4]), .ZN(n220) );
  OR2_X1 U391 ( .A1(B[0]), .A2(A[0]), .ZN(n475) );
  OAI211_X1 U392 ( .C1(A[1]), .C2(B[1]), .A(B[0]), .B(A[0]), .ZN(n474) );
  NAND2_X1 U393 ( .A1(B[1]), .A2(A[1]), .ZN(n317) );
  NAND2_X1 U394 ( .A1(B[5]), .A2(A[5]), .ZN(n103) );
  NAND2_X1 U395 ( .A1(B[4]), .A2(A[4]), .ZN(n151) );
  NAND2_X1 U396 ( .A1(B[6]), .A2(A[6]), .ZN(n96) );
  NAND2_X1 U397 ( .A1(B[2]), .A2(A[2]), .ZN(n257) );
  NAND4_X1 U398 ( .A1(n425), .A2(n90), .A3(n426), .A4(n427), .ZN(n416) );
  OR2_X1 U399 ( .A1(B[9]), .A2(A[9]), .ZN(n425) );
  NAND2_X1 U400 ( .A1(B[3]), .A2(A[3]), .ZN(n260) );
  NAND2_X1 U402 ( .A1(B[0]), .A2(A[0]), .ZN(n394) );
  OR2_X1 U403 ( .A1(B[11]), .A2(A[11]), .ZN(n427) );
  NAND2_X1 U404 ( .A1(B[7]), .A2(A[7]), .ZN(n99) );
  NAND2_X1 U405 ( .A1(B[13]), .A2(A[13]), .ZN(n436) );
  NOR2_X1 U406 ( .A1(A[13]), .A2(B[13]), .ZN(n434) );
  NAND2_X1 U407 ( .A1(net493832), .A2(n41), .ZN(net493830) );
  NOR2_X1 U408 ( .A1(n10), .A2(net493835), .ZN(n251) );
  NAND2_X1 U409 ( .A1(n449), .A2(n460), .ZN(n459) );
  AOI21_X1 U410 ( .B1(n228), .B2(n229), .A(n82), .ZN(n224) );
  NAND2_X1 U411 ( .A1(B[11]), .A2(A[11]), .ZN(n423) );
  OR2_X1 U412 ( .A1(B[11]), .A2(A[11]), .ZN(n451) );
  NAND2_X1 U413 ( .A1(n191), .A2(n192), .ZN(n168) );
  NAND2_X1 U414 ( .A1(net493866), .A2(net493865), .ZN(net493885) );
  NAND4_X1 U415 ( .A1(net493874), .A2(net493869), .A3(net493871), .A4(
        net493865), .ZN(net493809) );
  NAND2_X1 U416 ( .A1(n443), .A2(n435), .ZN(n441) );
  AND2_X1 U417 ( .A1(n443), .A2(n435), .ZN(n76) );
  NAND4_X1 U418 ( .A1(n22), .A2(n489), .A3(n351), .A4(n350), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n40), .B(net493850), .ZN(SUM[42]) );
  AND2_X1 U420 ( .A1(n222), .A2(n205), .ZN(n512) );
  NAND2_X1 U421 ( .A1(B[48]), .A2(A[48]), .ZN(n205) );
  AND2_X1 U422 ( .A1(n367), .A2(n358), .ZN(n3) );
  INV_X1 U423 ( .A(n358), .ZN(n539) );
  OAI21_X1 U424 ( .B1(n288), .B2(n23), .A(n290), .ZN(n279) );
  NAND2_X1 U425 ( .A1(n282), .A2(n283), .ZN(n280) );
  NAND2_X1 U426 ( .A1(n191), .A2(n516), .ZN(n513) );
  OR2_X1 U427 ( .A1(n515), .A2(n171), .ZN(n514) );
  INV_X1 U428 ( .A(n178), .ZN(n515) );
  AND2_X1 U429 ( .A1(n192), .A2(n178), .ZN(n516) );
  OR2_X1 U430 ( .A1(B[14]), .A2(A[14]), .ZN(n54) );
  NAND2_X1 U431 ( .A1(A[14]), .A2(B[14]), .ZN(n437) );
  OR2_X1 U432 ( .A1(A[14]), .A2(B[14]), .ZN(n432) );
  OAI21_X1 U433 ( .B1(n134), .B2(n530), .A(n136), .ZN(n132) );
  XNOR2_X1 U434 ( .A(n163), .B(n162), .ZN(SUM[56]) );
  OAI21_X1 U435 ( .B1(n554), .B2(n530), .A(n142), .ZN(n159) );
  INV_X1 U436 ( .A(n162), .ZN(n530) );
  XNOR2_X1 U437 ( .A(net538274), .B(net493856), .ZN(SUM[41]) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(SUM[23]) );
  OAI21_X1 U439 ( .B1(n523), .B2(n566), .A(net493872), .ZN(net537204) );
  NOR2_X1 U440 ( .A1(n86), .A2(n587), .ZN(n452) );
  NOR2_X1 U441 ( .A1(n586), .A2(n86), .ZN(n84) );
  OAI211_X1 U442 ( .C1(n86), .C2(n91), .A(n449), .B(n87), .ZN(n448) );
  OAI21_X1 U443 ( .B1(n83), .B2(n86), .A(n87), .ZN(n461) );
  AOI21_X1 U444 ( .B1(n289), .B2(n293), .A(n577), .ZN(n324) );
  AND2_X1 U445 ( .A1(n479), .A2(B[27]), .ZN(n11) );
  INV_X1 U446 ( .A(A[27]), .ZN(n574) );
  INV_X1 U447 ( .A(n267), .ZN(n569) );
  NAND2_X1 U448 ( .A1(B[19]), .A2(A[19]), .ZN(n382) );
  OR2_X1 U449 ( .A1(B[19]), .A2(A[19]), .ZN(n386) );
  NAND2_X1 U450 ( .A1(n164), .A2(n165), .ZN(n162) );
  INV_X1 U451 ( .A(n31), .ZN(n573) );
  AND3_X1 U452 ( .A1(n292), .A2(n71), .A3(n293), .ZN(n300) );
  XNOR2_X1 U453 ( .A(n71), .B(n407), .ZN(SUM[16]) );
  INV_X1 U454 ( .A(n71), .ZN(n521) );
  XNOR2_X1 U455 ( .A(n459), .B(n458), .ZN(SUM[11]) );
  NAND2_X1 U456 ( .A1(n19), .A2(n437), .ZN(n18) );
  NAND4_X1 U457 ( .A1(n279), .A2(n278), .A3(n280), .A4(n281), .ZN(n237) );
  AOI21_X1 U458 ( .B1(n201), .B2(n202), .A(n543), .ZN(n191) );
  INV_X1 U459 ( .A(net493790), .ZN(n557) );
  NAND2_X1 U460 ( .A1(n362), .A2(n336), .ZN(n368) );
  AND2_X1 U461 ( .A1(n362), .A2(n363), .ZN(n356) );
  NOR2_X1 U462 ( .A1(n542), .A2(n544), .ZN(n201) );
  NAND2_X1 U463 ( .A1(n183), .A2(n179), .ZN(n182) );
  NAND2_X1 U464 ( .A1(n331), .A2(n336), .ZN(n294) );
  NAND2_X1 U465 ( .A1(n249), .A2(n231), .ZN(n247) );
  OAI21_X1 U466 ( .B1(n517), .B2(n403), .A(n397), .ZN(n396) );
  INV_X1 U467 ( .A(n398), .ZN(n517) );
  XNOR2_X1 U468 ( .A(n396), .B(n395), .ZN(SUM[19]) );
  XNOR2_X1 U469 ( .A(n181), .B(n182), .ZN(SUM[55]) );
  XNOR2_X1 U470 ( .A(net493891), .B(net537204), .ZN(SUM[38]) );
  NAND2_X1 U471 ( .A1(n274), .A2(n271), .ZN(n66) );
  AOI21_X1 U472 ( .B1(n237), .B2(n272), .A(n568), .ZN(n75) );
  NAND2_X1 U473 ( .A1(n308), .A2(n392), .ZN(n406) );
  INV_X1 U474 ( .A(n415), .ZN(n534) );
  AND3_X1 U475 ( .A1(n432), .A2(n421), .A3(n415), .ZN(n419) );
  NAND2_X1 U476 ( .A1(n40), .A2(net493837), .ZN(n42) );
  NAND2_X1 U477 ( .A1(A[39]), .A2(B[39]), .ZN(net493866) );
  XNOR2_X1 U478 ( .A(n344), .B(n345), .ZN(SUM[27]) );
  NAND4_X1 U479 ( .A1(n490), .A2(n333), .A3(n334), .A4(n332), .ZN(n296) );
  NAND4_X1 U480 ( .A1(n333), .A2(n336), .A3(n332), .A4(n331), .ZN(n350) );
  INV_X1 U481 ( .A(n333), .ZN(n579) );
  OAI21_X1 U482 ( .B1(n323), .B2(n578), .A(n324), .ZN(n314) );
  NOR2_X1 U483 ( .A1(n307), .A2(n487), .ZN(n301) );
  OAI21_X1 U484 ( .B1(n521), .B2(n307), .A(n43), .ZN(n60) );
  NOR2_X1 U485 ( .A1(n483), .A2(B[18]), .ZN(n403) );
  OAI21_X1 U486 ( .B1(n521), .B2(n307), .A(n63), .ZN(n364) );
  NAND2_X1 U487 ( .A1(B[18]), .A2(n483), .ZN(n397) );
  OR2_X1 U488 ( .A1(B[18]), .A2(A[18]), .ZN(n384) );
  XNOR2_X1 U489 ( .A(n160), .B(n159), .ZN(SUM[57]) );
  INV_X1 U490 ( .A(n159), .ZN(n529) );
  NAND2_X1 U491 ( .A1(B[55]), .A2(A[55]), .ZN(n176) );
  OAI21_X1 U492 ( .B1(n531), .B2(n544), .A(n207), .ZN(n211) );
  XNOR2_X1 U493 ( .A(n462), .B(n461), .ZN(SUM[10]) );
  NAND2_X1 U494 ( .A1(n426), .A2(n461), .ZN(n460) );
  NAND2_X1 U495 ( .A1(B[8]), .A2(A[8]), .ZN(n91) );
  INV_X1 U496 ( .A(n35), .ZN(n524) );
  NAND2_X1 U497 ( .A1(A[33]), .A2(B[33]), .ZN(n270) );
  INV_X1 U498 ( .A(net493809), .ZN(n556) );
  XNOR2_X1 U499 ( .A(n444), .B(n445), .ZN(SUM[12]) );
  NAND2_X1 U500 ( .A1(n414), .A2(n444), .ZN(n443) );
  NAND2_X1 U501 ( .A1(n364), .A2(n367), .ZN(n376) );
  NAND2_X1 U502 ( .A1(net493824), .A2(n238), .ZN(n249) );
  OAI211_X1 U503 ( .C1(n533), .C2(n409), .A(n410), .B(n413), .ZN(n71) );
  OAI211_X1 U504 ( .C1(n533), .C2(n409), .A(n410), .B(n413), .ZN(n308) );
  INV_X1 U505 ( .A(n28), .ZN(n520) );
  NAND2_X1 U506 ( .A1(n28), .A2(n287), .ZN(n24) );
  AOI21_X1 U507 ( .B1(n292), .B2(n314), .A(n582), .ZN(n28) );
  OR2_X1 U508 ( .A1(B[25]), .A2(A[25]), .ZN(n340) );
  NAND2_X1 U509 ( .A1(A[25]), .A2(B[25]), .ZN(n341) );
  AND4_X1 U510 ( .A1(n381), .A2(n380), .A3(n379), .A4(n382), .ZN(n43) );
  AND4_X1 U511 ( .A1(n380), .A2(n381), .A3(n379), .A4(n382), .ZN(n63) );
  AOI21_X1 U512 ( .B1(n485), .B2(n556), .A(n557), .ZN(n227) );
  XNOR2_X1 U513 ( .A(n50), .B(n275), .ZN(SUM[34]) );
  NAND2_X1 U514 ( .A1(n50), .A2(n265), .ZN(n274) );
  INV_X1 U516 ( .A(n75), .ZN(n532) );
  OAI21_X1 U517 ( .B1(n75), .B2(n571), .A(n270), .ZN(n50) );
  XNOR2_X1 U518 ( .A(n210), .B(n211), .ZN(SUM[51]) );
  NAND4_X1 U519 ( .A1(n556), .A2(net538113), .A3(n560), .A4(n39), .ZN(
        net493779) );
  NAND4_X1 U520 ( .A1(n386), .A2(n384), .A3(n385), .A4(n492), .ZN(n381) );
  XNOR2_X1 U521 ( .A(n347), .B(n349), .ZN(SUM[26]) );
  AOI21_X1 U522 ( .B1(n334), .B2(n347), .A(n576), .ZN(n344) );
  NAND2_X1 U523 ( .A1(n294), .A2(n330), .ZN(n354) );
  INV_X1 U524 ( .A(n330), .ZN(n518) );
  NAND2_X1 U525 ( .A1(A[23]), .A2(B[23]), .ZN(n362) );
  INV_X1 U526 ( .A(A[23]), .ZN(n572) );
  XNOR2_X1 U527 ( .A(n439), .B(n440), .ZN(SUM[14]) );
  NAND2_X1 U528 ( .A1(n439), .A2(n54), .ZN(n19) );
  NAND2_X1 U529 ( .A1(n447), .A2(n448), .ZN(n2) );
  NAND2_X1 U530 ( .A1(n447), .A2(n448), .ZN(n422) );
  NAND2_X1 U531 ( .A1(A[10]), .A2(B[10]), .ZN(n449) );
  XNOR2_X1 U532 ( .A(net493858), .B(net493861), .ZN(SUM[40]) );
  OAI21_X1 U534 ( .B1(n34), .B2(n565), .A(net493839), .ZN(n40) );
  INV_X1 U535 ( .A(n488), .ZN(n522) );
  NAND2_X1 U536 ( .A1(n204), .A2(n197), .ZN(n210) );
  AND3_X1 U537 ( .A1(n195), .A2(n196), .A3(n197), .ZN(n194) );
  INV_X1 U538 ( .A(n197), .ZN(n542) );
  INV_X1 U539 ( .A(net493785), .ZN(n560) );
  OAI21_X1 U540 ( .B1(n227), .B2(net493785), .A(net493786), .ZN(n226) );
  OAI21_X1 U541 ( .B1(n522), .B2(net493785), .A(net493786), .ZN(net493824) );
  INV_X1 U542 ( .A(net493791), .ZN(n561) );
  NOR2_X1 U543 ( .A1(net493791), .A2(net493805), .ZN(n39) );
  AND2_X1 U544 ( .A1(A[47]), .A2(B[47]), .ZN(n82) );
  INV_X1 U545 ( .A(net493900), .ZN(n523) );
  AOI21_X1 U546 ( .B1(net493900), .B2(net493869), .A(n567), .ZN(n35) );
  OAI21_X1 U547 ( .B1(n16), .B2(n555), .A(net493873), .ZN(net493900) );
  NAND4_X1 U548 ( .A1(n266), .A2(n273), .A3(n265), .A4(n272), .ZN(net493805)
         );
  NAND2_X1 U549 ( .A1(n265), .A2(n266), .ZN(n263) );
  XNOR2_X1 U550 ( .A(net493845), .B(n252), .ZN(SUM[43]) );
  NAND2_X1 U551 ( .A1(n42), .A2(n41), .ZN(net493845) );
  OAI21_X1 U552 ( .B1(n9), .B2(net493864), .A(net493865), .ZN(net493790) );
  NAND2_X1 U553 ( .A1(net493866), .A2(net493867), .ZN(net493864) );
  AOI21_X1 U554 ( .B1(net493841), .B2(net493858), .A(n558), .ZN(n34) );
  OAI21_X1 U555 ( .B1(n497), .B2(net493809), .A(net493790), .ZN(net493858) );
  NAND2_X1 U557 ( .A1(n169), .A2(n184), .ZN(n183) );
  NAND2_X1 U558 ( .A1(net493832), .A2(net493831), .ZN(n252) );
  NAND4_X1 U559 ( .A1(net493841), .A2(net493836), .A3(net493837), .A4(
        net493831), .ZN(net493785) );
  NAND2_X1 U560 ( .A1(B[43]), .A2(A[43]), .ZN(net493832) );
  INV_X1 U561 ( .A(n213), .ZN(n531) );
  NAND2_X1 U562 ( .A1(n193), .A2(n194), .ZN(n192) );
  XNOR2_X1 U564 ( .A(n193), .B(n223), .ZN(SUM[48]) );
  NAND2_X1 U565 ( .A1(n193), .A2(n200), .ZN(n222) );
  XNOR2_X1 U566 ( .A(n241), .B(n242), .ZN(SUM[47]) );
  AOI21_X1 U569 ( .B1(n236), .B2(n243), .A(n563), .ZN(n241) );
  OAI21_X1 U570 ( .B1(n251), .B2(net493830), .A(net493831), .ZN(net493786) );
endmodule


module RCA_NBIT64_12 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_12_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), 
        .SUM({Co, S}) );
endmodule


module RCA_NBIT64_11_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net494959, net494954, net494951, net494949, net494943, net494942,
         net494937, net494936, net494931, net494930, net494915, net494900,
         net494899, net494888, net494882, net494881, net494879, net494878,
         net494876, net535402, net537213, net537812, net537811, net494929,
         net494895, net494955, net494945, net494939, net494902, net494938,
         net494935, net494933, net538681, net494958, net494944, net494934,
         net494928, net494892, net494884, net494883, net494922, net494921,
         net494917, net494911, net494904, net494903, net494894, net494893, n3,
         n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n17, n18, n21, n24,
         n25, n27, n29, n30, n37, n39, n40, n41, n45, n47, n48, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n63, n64, n66, n67, n68, n70,
         n71, n72, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n110, n111, n112, n113,
         n115, n116, n117, n118, n119, n120, n122, n123, n126, n127, n129,
         n130, n131, n133, n134, n135, n136, n138, n139, n141, n142, n143,
         n145, n146, n147, n150, n151, n152, n153, n154, n156, n157, n158,
         n159, n160, n162, n164, n166, n168, n170, n171, n172, n173, n174,
         n175, n177, n178, n179, n182, n183, n184, n185, n186, n187, n188,
         n192, n194, n196, n198, n199, n200, n202, n204, n205, n206, n207,
         n208, n209, n210, n212, n213, n214, n217, n218, n220, n221, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n243, n244, n245, n246, n247,
         n248, n249, n252, n254, n256, n257, n258, n259, n261, n262, n263,
         n264, n265, n266, n267, n269, n270, n271, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n284, n285, n286, n288, n289,
         n290, n292, n294, n295, n296, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n313, n314, n315,
         n317, n318, n319, n320, n321, n322, n324, n325, n326, n328, n329,
         n330, n331, n336, n337, n339, n340, n341, n342, n343, n344, n347,
         n348, n349, n353, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n373, n374, n376, n377,
         n378, n380, n381, n382, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n411, n412, n413, n414, n415, n416, n417,
         n419, n421, n423, n424, n425, n426, n427, n429, n430, n431, n433,
         n434, n435, n436, n438, n439, n440, n441, n442, n443, n444, n445,
         n448, n449, n450, n452, n453, n455, n456, n457, n459, n460, n461,
         n462, n464, n465, n466, n467, n468, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596;

  OR2_X2 U18 ( .A1(A[43]), .A2(B[43]), .ZN(net494929) );
  OR2_X2 U109 ( .A1(A[42]), .A2(B[42]), .ZN(net494935) );
  NAND3_X1 U134 ( .A1(n259), .A2(n258), .A3(n14), .ZN(n225) );
  OR2_X2 U136 ( .A1(B[34]), .A2(A[34]), .ZN(n258) );
  OR2_X2 U360 ( .A1(A[22]), .A2(B[22]), .ZN(n359) );
  NAND3_X1 U559 ( .A1(n273), .A2(n275), .A3(n274), .ZN(n226) );
  NAND3_X1 U561 ( .A1(n84), .A2(n303), .A3(n304), .ZN(n282) );
  NAND3_X1 U588 ( .A1(n86), .A2(n96), .A3(n426), .ZN(n438) );
  NAND3_X1 U589 ( .A1(n449), .A2(n448), .A3(n450), .ZN(n442) );
  OR2_X2 U19 ( .A1(B[13]), .A2(A[13]), .ZN(n415) );
  OR2_X2 U30 ( .A1(A[41]), .A2(B[41]), .ZN(net494933) );
  OR2_X2 U77 ( .A1(B[46]), .A2(A[46]), .ZN(net494894) );
  OR2_X2 U325 ( .A1(A[19]), .A2(B[19]), .ZN(n382) );
  OR2_X2 U330 ( .A1(B[18]), .A2(A[18]), .ZN(n381) );
  OR2_X2 U332 ( .A1(B[54]), .A2(A[54]), .ZN(n182) );
  OR2_X2 U346 ( .A1(B[37]), .A2(A[37]), .ZN(n233) );
  OR2_X2 U380 ( .A1(A[12]), .A2(B[12]), .ZN(n440) );
  CLKBUF_X1 U2 ( .A(n288), .Z(n472) );
  OR2_X1 U3 ( .A1(B[21]), .A2(A[21]), .ZN(n360) );
  OR2_X1 U4 ( .A1(B[20]), .A2(A[20]), .ZN(n365) );
  OR2_X1 U5 ( .A1(B[24]), .A2(A[24]), .ZN(n336) );
  OR2_X1 U6 ( .A1(B[28]), .A2(A[28]), .ZN(n300) );
  OR2_X1 U7 ( .A1(B[29]), .A2(A[29]), .ZN(n301) );
  AND2_X1 U8 ( .A1(n464), .A2(n392), .ZN(SUM[0]) );
  OR2_X1 U9 ( .A1(B[40]), .A2(A[40]), .ZN(net494938) );
  OR2_X1 U10 ( .A1(B[32]), .A2(A[32]), .ZN(n256) );
  OR2_X1 U11 ( .A1(B[36]), .A2(A[36]), .ZN(n238) );
  OR2_X1 U12 ( .A1(A[39]), .A2(B[39]), .ZN(n229) );
  OR2_X1 U13 ( .A1(B[45]), .A2(A[45]), .ZN(net494893) );
  OR2_X1 U14 ( .A1(B[44]), .A2(A[44]), .ZN(net494892) );
  OR2_X1 U15 ( .A1(B[48]), .A2(A[48]), .ZN(n221) );
  NOR2_X1 U16 ( .A1(A[49]), .A2(B[49]), .ZN(n87) );
  OR2_X1 U17 ( .A1(B[50]), .A2(A[50]), .ZN(n204) );
  OR2_X1 U20 ( .A1(B[53]), .A2(A[53]), .ZN(n184) );
  OR2_X1 U21 ( .A1(B[52]), .A2(A[52]), .ZN(n183) );
  OR2_X1 U22 ( .A1(B[58]), .A2(A[58]), .ZN(n150) );
  CLKBUF_X1 U23 ( .A(n27), .Z(n473) );
  AND2_X1 U24 ( .A1(n202), .A2(n526), .ZN(n474) );
  AND2_X1 U25 ( .A1(n17), .A2(n13), .ZN(n475) );
  BUF_X1 U26 ( .A(A[11]), .Z(n476) );
  INV_X1 U27 ( .A(n555), .ZN(n477) );
  OAI221_X1 U28 ( .B1(n29), .B2(n225), .C1(n261), .C2(n560), .A(n262), .ZN(
        n478) );
  OAI221_X1 U29 ( .B1(n29), .B2(n225), .C1(n261), .C2(n560), .A(n262), .ZN(
        n479) );
  OAI221_X1 U31 ( .B1(n29), .B2(n225), .C1(n261), .C2(n560), .A(n262), .ZN(
        n237) );
  NAND2_X1 U32 ( .A1(n3), .A2(n475), .ZN(n273) );
  OR2_X1 U33 ( .A1(A[11]), .A2(B[11]), .ZN(n450) );
  NOR2_X1 U34 ( .A1(B[27]), .A2(A[27]), .ZN(n85) );
  OR2_X1 U35 ( .A1(n276), .A2(n277), .ZN(n480) );
  NAND2_X1 U36 ( .A1(n480), .A2(n82), .ZN(n275) );
  CLKBUF_X1 U37 ( .A(n342), .Z(n481) );
  OR2_X1 U38 ( .A1(B[30]), .A2(A[30]), .ZN(n482) );
  OR2_X1 U39 ( .A1(B[30]), .A2(A[30]), .ZN(n483) );
  OR2_X1 U40 ( .A1(B[30]), .A2(A[30]), .ZN(n302) );
  NAND3_X1 U41 ( .A1(n449), .A2(n448), .A3(n450), .ZN(n484) );
  NAND2_X1 U42 ( .A1(n385), .A2(n386), .ZN(n485) );
  XNOR2_X1 U43 ( .A(n344), .B(n486), .ZN(SUM[27]) );
  NOR2_X1 U44 ( .A1(n542), .A2(n85), .ZN(n486) );
  AND2_X1 U45 ( .A1(A[15]), .A2(B[15]), .ZN(n487) );
  NAND4_X2 U46 ( .A1(n382), .A2(n380), .A3(n381), .A4(n399), .ZN(n306) );
  XNOR2_X1 U47 ( .A(n488), .B(n431), .ZN(SUM[15]) );
  AND2_X1 U48 ( .A1(n61), .A2(n60), .ZN(n488) );
  AND2_X1 U49 ( .A1(net494921), .A2(net494902), .ZN(n489) );
  XNOR2_X1 U50 ( .A(n267), .B(n490), .ZN(SUM[35]) );
  NAND2_X1 U51 ( .A1(n262), .A2(n18), .ZN(n490) );
  OR2_X1 U52 ( .A1(n405), .A2(n24), .ZN(n491) );
  NAND2_X1 U53 ( .A1(n491), .A2(n407), .ZN(n52) );
  OR2_X1 U54 ( .A1(A[31]), .A2(B[31]), .ZN(n492) );
  OR2_X1 U55 ( .A1(A[31]), .A2(B[31]), .ZN(n298) );
  AND2_X1 U56 ( .A1(n294), .A2(n295), .ZN(n493) );
  AND2_X1 U57 ( .A1(n317), .A2(n493), .ZN(n310) );
  XNOR2_X1 U58 ( .A(net537213), .B(n494), .ZN(SUM[42]) );
  NAND2_X1 U59 ( .A1(net494935), .A2(net494931), .ZN(n494) );
  NAND2_X1 U60 ( .A1(n83), .A2(n479), .ZN(n495) );
  AND2_X1 U61 ( .A1(n204), .A2(n205), .ZN(n496) );
  AOI21_X1 U62 ( .B1(n331), .B2(n336), .A(n543), .ZN(n497) );
  AOI21_X1 U63 ( .B1(n331), .B2(n336), .A(n543), .ZN(n77) );
  AND3_X1 U64 ( .A1(n198), .A2(n199), .A3(n200), .ZN(n498) );
  AND3_X1 U65 ( .A1(n198), .A2(n199), .A3(n200), .ZN(n172) );
  OR2_X1 U66 ( .A1(B[38]), .A2(A[38]), .ZN(n499) );
  OR2_X1 U67 ( .A1(A[38]), .A2(B[38]), .ZN(n234) );
  XNOR2_X1 U68 ( .A(n500), .B(n212), .ZN(SUM[51]) );
  NAND2_X1 U69 ( .A1(n205), .A2(n199), .ZN(n500) );
  OAI21_X1 U70 ( .B1(n497), .B2(n544), .A(n481), .ZN(n501) );
  XNOR2_X1 U71 ( .A(n48), .B(n502), .ZN(SUM[23]) );
  AND2_X1 U72 ( .A1(n64), .A2(n364), .ZN(n502) );
  XNOR2_X1 U73 ( .A(n503), .B(n252), .ZN(SUM[37]) );
  NAND2_X1 U74 ( .A1(n233), .A2(n235), .ZN(n503) );
  NAND2_X1 U75 ( .A1(n496), .A2(n474), .ZN(n200) );
  XOR2_X1 U76 ( .A(n504), .B(n45), .Z(SUM[13]) );
  AND2_X1 U78 ( .A1(n415), .A2(n416), .ZN(n504) );
  XNOR2_X1 U79 ( .A(n505), .B(n188), .ZN(SUM[54]) );
  NAND2_X1 U80 ( .A1(n182), .A2(n179), .ZN(n505) );
  XOR2_X1 U81 ( .A(n54), .B(n506), .Z(SUM[38]) );
  AND2_X1 U82 ( .A1(n499), .A2(n231), .ZN(n506) );
  XOR2_X1 U83 ( .A(n507), .B(n214), .Z(SUM[50]) );
  AND2_X1 U84 ( .A1(n204), .A2(n209), .ZN(n507) );
  XOR2_X1 U85 ( .A(n508), .B(n526), .Z(SUM[48]) );
  AND2_X1 U86 ( .A1(n221), .A2(n208), .ZN(n508) );
  XOR2_X1 U87 ( .A(n29), .B(n509), .Z(SUM[32]) );
  NAND2_X1 U88 ( .A1(n264), .A2(n256), .ZN(n509) );
  XOR2_X1 U89 ( .A(n510), .B(net494917), .Z(SUM[45]) );
  AND2_X1 U90 ( .A1(net494893), .A2(net494903), .ZN(n510) );
  XOR2_X1 U91 ( .A(n517), .B(n511), .Z(SUM[18]) );
  NAND2_X1 U92 ( .A1(n381), .A2(n389), .ZN(n511) );
  XOR2_X1 U93 ( .A(n512), .B(net537811), .Z(SUM[44]) );
  AND2_X1 U94 ( .A1(net494892), .A2(net494902), .ZN(n512) );
  AND4_X2 U95 ( .A1(n229), .A2(n233), .A3(n499), .A4(n238), .ZN(n83) );
  OR2_X1 U96 ( .A1(B[26]), .A2(A[26]), .ZN(n303) );
  XOR2_X1 U97 ( .A(n453), .B(n513), .Z(SUM[11]) );
  AND2_X1 U98 ( .A1(n452), .A2(n455), .ZN(n513) );
  AOI21_X1 U99 ( .B1(n289), .B2(n290), .A(n548), .ZN(n41) );
  OAI21_X1 U100 ( .B1(n421), .B2(n581), .A(n423), .ZN(n24) );
  INV_X1 U101 ( .A(n53), .ZN(n528) );
  AOI21_X1 U102 ( .B1(n289), .B2(n290), .A(n548), .ZN(n274) );
  OAI21_X1 U103 ( .B1(n421), .B2(n581), .A(n423), .ZN(n406) );
  NOR2_X1 U104 ( .A1(n528), .A2(n306), .ZN(n299) );
  AND3_X1 U105 ( .A1(n273), .A2(n41), .A3(n275), .ZN(n29) );
  INV_X1 U106 ( .A(n305), .ZN(n536) );
  INV_X1 U107 ( .A(n4), .ZN(n581) );
  INV_X1 U108 ( .A(n30), .ZN(n526) );
  NAND2_X1 U110 ( .A1(n71), .A2(n72), .ZN(n55) );
  OAI21_X1 U111 ( .B1(n592), .B2(n430), .A(n429), .ZN(n96) );
  NOR2_X1 U112 ( .A1(n425), .A2(n419), .ZN(n421) );
  NAND2_X1 U113 ( .A1(n86), .A2(n426), .ZN(n419) );
  AOI21_X1 U114 ( .B1(n586), .B2(n427), .A(n585), .ZN(n425) );
  INV_X1 U115 ( .A(n429), .ZN(n585) );
  INV_X1 U116 ( .A(n427), .ZN(n592) );
  INV_X1 U117 ( .A(n430), .ZN(n586) );
  NOR2_X1 U118 ( .A1(n113), .A2(n568), .ZN(SUM[64]) );
  NAND2_X1 U119 ( .A1(n365), .A2(n361), .ZN(n376) );
  NAND2_X1 U120 ( .A1(n258), .A2(n266), .ZN(n271) );
  NAND2_X1 U121 ( .A1(n348), .A2(n303), .ZN(n349) );
  XNOR2_X1 U122 ( .A(n373), .B(n374), .ZN(SUM[21]) );
  NOR2_X1 U123 ( .A1(n537), .A2(n535), .ZN(n374) );
  INV_X1 U124 ( .A(n363), .ZN(n537) );
  INV_X1 U125 ( .A(n233), .ZN(n558) );
  INV_X1 U126 ( .A(n236), .ZN(n552) );
  NAND2_X1 U127 ( .A1(n230), .A2(n231), .ZN(n228) );
  NOR2_X1 U128 ( .A1(n12), .A2(n232), .ZN(n227) );
  AND2_X1 U129 ( .A1(n235), .A2(n236), .ZN(n12) );
  NAND2_X1 U130 ( .A1(n292), .A2(n492), .ZN(n308) );
  NAND2_X1 U131 ( .A1(n301), .A2(n302), .ZN(n311) );
  NAND2_X1 U132 ( .A1(net494938), .A2(net494937), .ZN(net494958) );
  AND2_X1 U133 ( .A1(n265), .A2(n257), .ZN(n7) );
  XOR2_X1 U135 ( .A(n514), .B(n478), .Z(SUM[36]) );
  AND2_X1 U137 ( .A1(n238), .A2(n236), .ZN(n514) );
  NAND2_X1 U138 ( .A1(n133), .A2(n122), .ZN(n135) );
  NAND2_X1 U139 ( .A1(n129), .A2(n120), .ZN(n131) );
  NAND2_X1 U140 ( .A1(n300), .A2(n294), .ZN(n328) );
  NAND2_X1 U141 ( .A1(n359), .A2(n362), .ZN(n368) );
  NOR2_X1 U142 ( .A1(n547), .A2(n546), .ZN(n315) );
  AOI21_X1 U143 ( .B1(n313), .B2(n301), .A(n550), .ZN(n314) );
  INV_X1 U144 ( .A(n296), .ZN(n547) );
  XNOR2_X1 U145 ( .A(n53), .B(n404), .ZN(SUM[16]) );
  NAND2_X1 U146 ( .A1(n401), .A2(n380), .ZN(n404) );
  OAI211_X1 U147 ( .C1(n580), .C2(n438), .A(n439), .B(n417), .ZN(n45) );
  XNOR2_X1 U148 ( .A(n325), .B(n326), .ZN(SUM[29]) );
  NOR2_X1 U149 ( .A1(n550), .A2(n549), .ZN(n326) );
  INV_X1 U150 ( .A(n294), .ZN(n545) );
  OAI211_X1 U151 ( .C1(n549), .C2(n294), .A(n295), .B(n296), .ZN(n290) );
  NAND2_X1 U152 ( .A1(n382), .A2(n286), .ZN(n393) );
  OAI21_X1 U153 ( .B1(n55), .B2(n533), .A(n389), .ZN(n394) );
  INV_X1 U154 ( .A(n381), .ZN(n533) );
  NOR2_X1 U155 ( .A1(n579), .A2(n87), .ZN(n218) );
  INV_X1 U156 ( .A(n147), .ZN(n572) );
  NAND2_X1 U157 ( .A1(n424), .A2(n413), .ZN(n434) );
  NAND2_X1 U158 ( .A1(n67), .A2(n68), .ZN(n48) );
  OR2_X1 U159 ( .A1(n539), .A2(n359), .ZN(n68) );
  INV_X1 U160 ( .A(n279), .ZN(n542) );
  AOI21_X1 U161 ( .B1(n83), .B2(n223), .A(n553), .ZN(net494882) );
  OAI21_X1 U162 ( .B1(n560), .B2(n261), .A(n262), .ZN(n223) );
  OAI21_X1 U163 ( .B1(n520), .B2(n576), .A(n146), .ZN(n160) );
  OAI21_X1 U164 ( .B1(n527), .B2(n87), .A(n210), .ZN(n214) );
  NOR2_X1 U165 ( .A1(n575), .A2(n576), .ZN(n164) );
  INV_X1 U166 ( .A(n146), .ZN(n575) );
  INV_X1 U167 ( .A(n179), .ZN(n565) );
  XOR2_X1 U168 ( .A(n51), .B(n515), .Z(SUM[24]) );
  AND2_X1 U169 ( .A1(n353), .A2(n336), .ZN(n515) );
  AOI21_X1 U170 ( .B1(net494939), .B2(net494938), .A(n557), .ZN(net494949) );
  XNOR2_X1 U171 ( .A(net494951), .B(net494954), .ZN(SUM[41]) );
  NAND2_X1 U172 ( .A1(net494955), .A2(net494937), .ZN(net494951) );
  XNOR2_X1 U173 ( .A(n77), .B(n516), .ZN(SUM[25]) );
  AND2_X1 U174 ( .A1(n342), .A2(n337), .ZN(n516) );
  XNOR2_X1 U175 ( .A(net494915), .B(net537812), .ZN(SUM[46]) );
  NAND2_X1 U176 ( .A1(net494894), .A2(net494904), .ZN(net494915) );
  XNOR2_X1 U177 ( .A(n162), .B(n160), .ZN(SUM[58]) );
  NAND2_X1 U178 ( .A1(n150), .A2(n147), .ZN(n162) );
  XNOR2_X1 U179 ( .A(n444), .B(n445), .ZN(SUM[12]) );
  NAND2_X1 U180 ( .A1(n440), .A2(n417), .ZN(n444) );
  NAND2_X1 U181 ( .A1(n4), .A2(n438), .ZN(n445) );
  NAND2_X1 U182 ( .A1(n71), .A2(n72), .ZN(n517) );
  XNOR2_X1 U183 ( .A(n524), .B(n168), .ZN(SUM[56]) );
  NOR2_X1 U184 ( .A1(n577), .A2(n578), .ZN(n168) );
  INV_X1 U185 ( .A(n145), .ZN(n577) );
  INV_X1 U186 ( .A(n150), .ZN(n573) );
  NAND4_X1 U187 ( .A1(n64), .A2(n360), .A3(n359), .A4(n365), .ZN(n305) );
  NAND2_X1 U188 ( .A1(n269), .A2(n266), .ZN(n267) );
  AOI21_X1 U189 ( .B1(n280), .B2(n281), .A(n282), .ZN(n276) );
  NAND2_X1 U190 ( .A1(n278), .A2(n279), .ZN(n277) );
  AND3_X1 U191 ( .A1(n298), .A2(n302), .A3(n58), .ZN(n82) );
  OAI21_X1 U192 ( .B1(n523), .B2(n88), .A(n123), .ZN(n134) );
  OAI21_X1 U193 ( .B1(n522), .B2(n570), .A(n122), .ZN(n130) );
  OAI211_X1 U194 ( .C1(n576), .C2(n145), .A(n146), .B(n147), .ZN(n143) );
  OAI211_X1 U195 ( .C1(n556), .C2(net494902), .A(net494903), .B(net494904), 
        .ZN(net494900) );
  INV_X1 U196 ( .A(n353), .ZN(n543) );
  XNOR2_X1 U197 ( .A(n523), .B(n136), .ZN(SUM[60]) );
  NOR2_X1 U198 ( .A1(n571), .A2(n88), .ZN(n136) );
  INV_X1 U199 ( .A(n123), .ZN(n571) );
  XNOR2_X1 U200 ( .A(n126), .B(n127), .ZN(SUM[63]) );
  NAND2_X1 U201 ( .A1(n119), .A2(n115), .ZN(n126) );
  OAI21_X1 U202 ( .B1(n521), .B2(n569), .A(n120), .ZN(n127) );
  XNOR2_X1 U203 ( .A(n248), .B(n247), .ZN(SUM[39]) );
  NAND2_X1 U204 ( .A1(n249), .A2(n231), .ZN(n248) );
  OAI211_X1 U205 ( .C1(n583), .C2(n98), .A(n94), .B(n452), .ZN(n449) );
  XNOR2_X1 U206 ( .A(net494943), .B(net494942), .ZN(SUM[43]) );
  NAND2_X1 U207 ( .A1(net494930), .A2(net494929), .ZN(net494942) );
  NAND2_X1 U208 ( .A1(net494944), .A2(net494931), .ZN(net494943) );
  OAI21_X1 U209 ( .B1(n10), .B2(net494928), .A(net494929), .ZN(n21) );
  AND2_X1 U210 ( .A1(n536), .A2(n299), .ZN(n13) );
  AND3_X1 U211 ( .A1(n84), .A2(n303), .A3(n304), .ZN(n17) );
  AND3_X1 U212 ( .A1(n492), .A2(n482), .A3(n58), .ZN(n3) );
  AOI21_X1 U213 ( .B1(net494939), .B2(net494938), .A(n557), .ZN(n25) );
  OAI211_X1 U214 ( .C1(n567), .C2(n177), .A(n178), .B(n179), .ZN(n175) );
  NOR2_X1 U215 ( .A1(n288), .A2(n538), .ZN(n355) );
  OAI21_X1 U216 ( .B1(n578), .B2(n524), .A(n145), .ZN(n166) );
  INV_X1 U217 ( .A(n138), .ZN(n523) );
  AOI21_X1 U218 ( .B1(n142), .B2(n143), .A(n90), .ZN(n141) );
  NOR2_X1 U219 ( .A1(n538), .A2(n472), .ZN(n280) );
  INV_X1 U220 ( .A(n152), .ZN(n576) );
  NAND2_X1 U221 ( .A1(n11), .A2(net494929), .ZN(net494883) );
  AND3_X1 U222 ( .A1(net494935), .A2(net494933), .A3(net494938), .ZN(n11) );
  NAND2_X1 U223 ( .A1(n541), .A2(n590), .ZN(n304) );
  INV_X1 U224 ( .A(n170), .ZN(n524) );
  OAI211_X1 U225 ( .C1(n580), .C2(n438), .A(n439), .B(n417), .ZN(n436) );
  NOR2_X1 U226 ( .A1(n566), .A2(n567), .ZN(n192) );
  INV_X1 U227 ( .A(n178), .ZN(n566) );
  NOR2_X1 U228 ( .A1(n562), .A2(n563), .ZN(n196) );
  INV_X1 U229 ( .A(n177), .ZN(n562) );
  NAND2_X1 U230 ( .A1(net494899), .A2(net494900), .ZN(net494876) );
  NAND2_X1 U231 ( .A1(net535402), .A2(net494881), .ZN(net494879) );
  NAND2_X1 U232 ( .A1(n329), .A2(n330), .ZN(n318) );
  NAND4_X1 U233 ( .A1(n84), .A2(n303), .A3(n304), .A4(n51), .ZN(n330) );
  AND2_X1 U234 ( .A1(n278), .A2(n279), .ZN(n329) );
  AND4_X1 U235 ( .A1(net494895), .A2(net494893), .A3(net494894), .A4(net494892), .ZN(net535402) );
  INV_X1 U236 ( .A(n361), .ZN(n551) );
  NAND2_X1 U237 ( .A1(net494921), .A2(net494902), .ZN(net494917) );
  NAND2_X1 U238 ( .A1(n440), .A2(n441), .ZN(n439) );
  NAND2_X1 U239 ( .A1(n442), .A2(n443), .ZN(n441) );
  OAI21_X1 U240 ( .B1(n87), .B2(n208), .A(n209), .ZN(n206) );
  INV_X1 U241 ( .A(n184), .ZN(n567) );
  AND2_X1 U242 ( .A1(n363), .A2(n362), .ZN(n70) );
  NOR2_X1 U243 ( .A1(n87), .A2(n561), .ZN(n202) );
  NOR2_X1 U244 ( .A1(n75), .A2(n225), .ZN(n224) );
  AND3_X1 U245 ( .A1(net494933), .A2(net494934), .A3(net494935), .ZN(n10) );
  AND2_X1 U246 ( .A1(n484), .A2(n443), .ZN(n4) );
  AND2_X1 U247 ( .A1(n424), .A2(n76), .ZN(n423) );
  AND2_X1 U248 ( .A1(n415), .A2(n440), .ZN(n76) );
  AND2_X1 U249 ( .A1(n298), .A2(n483), .ZN(n289) );
  INV_X1 U250 ( .A(n364), .ZN(n538) );
  NAND2_X1 U251 ( .A1(n18), .A2(n258), .ZN(n261) );
  INV_X1 U252 ( .A(net494937), .ZN(n557) );
  NAND2_X1 U253 ( .A1(n400), .A2(n74), .ZN(n71) );
  AND2_X1 U254 ( .A1(n401), .A2(n398), .ZN(n74) );
  INV_X1 U255 ( .A(n292), .ZN(n548) );
  INV_X1 U256 ( .A(net494893), .ZN(n556) );
  INV_X1 U257 ( .A(n295), .ZN(n550) );
  INV_X1 U258 ( .A(n133), .ZN(n570) );
  INV_X1 U259 ( .A(n301), .ZN(n549) );
  INV_X1 U260 ( .A(n129), .ZN(n569) );
  INV_X1 U261 ( .A(n151), .ZN(n578) );
  XNOR2_X1 U262 ( .A(n5), .B(n6), .ZN(SUM[47]) );
  NAND2_X1 U263 ( .A1(net494904), .A2(net494911), .ZN(n5) );
  NAND2_X1 U264 ( .A1(n536), .A2(n284), .ZN(n281) );
  NAND2_X1 U265 ( .A1(n233), .A2(n234), .ZN(n232) );
  OR2_X1 U266 ( .A1(n532), .A2(n399), .ZN(n72) );
  INV_X1 U267 ( .A(n398), .ZN(n532) );
  INV_X1 U268 ( .A(n263), .ZN(n560) );
  OAI211_X1 U269 ( .C1(n78), .C2(n264), .A(n265), .B(n266), .ZN(n263) );
  AND2_X1 U270 ( .A1(n416), .A2(n413), .ZN(n63) );
  INV_X1 U271 ( .A(n210), .ZN(n579) );
  INV_X1 U272 ( .A(n221), .ZN(n561) );
  INV_X1 U273 ( .A(n183), .ZN(n563) );
  INV_X1 U274 ( .A(n348), .ZN(n540) );
  AND2_X1 U275 ( .A1(n301), .A2(n300), .ZN(n58) );
  AND2_X1 U276 ( .A1(n377), .A2(n378), .ZN(n79) );
  NAND2_X1 U277 ( .A1(n531), .A2(n53), .ZN(n378) );
  INV_X1 U278 ( .A(n306), .ZN(n531) );
  INV_X1 U279 ( .A(n264), .ZN(n559) );
  INV_X1 U280 ( .A(n482), .ZN(n546) );
  INV_X1 U281 ( .A(net494933), .ZN(n554) );
  INV_X1 U282 ( .A(n360), .ZN(n535) );
  INV_X1 U283 ( .A(n413), .ZN(n530) );
  INV_X1 U284 ( .A(n362), .ZN(n539) );
  XNOR2_X1 U285 ( .A(n99), .B(n100), .ZN(SUM[7]) );
  NAND2_X1 U286 ( .A1(n103), .A2(n104), .ZN(n99) );
  NAND2_X1 U287 ( .A1(n101), .A2(n102), .ZN(n100) );
  NAND2_X1 U288 ( .A1(n105), .A2(n106), .ZN(n104) );
  XNOR2_X1 U289 ( .A(n239), .B(n240), .ZN(SUM[3]) );
  OAI21_X1 U290 ( .B1(n595), .B2(n593), .A(n243), .ZN(n240) );
  NAND2_X1 U291 ( .A1(n245), .A2(n246), .ZN(n239) );
  INV_X1 U292 ( .A(n244), .ZN(n595) );
  XNOR2_X1 U293 ( .A(n91), .B(n92), .ZN(SUM[9]) );
  NAND2_X1 U294 ( .A1(n93), .A2(n94), .ZN(n91) );
  XNOR2_X1 U295 ( .A(n95), .B(n96), .ZN(SUM[8]) );
  NAND2_X1 U296 ( .A1(n97), .A2(n98), .ZN(n95) );
  XNOR2_X1 U297 ( .A(n217), .B(n427), .ZN(SUM[4]) );
  NAND2_X1 U298 ( .A1(n157), .A2(n156), .ZN(n217) );
  XNOR2_X1 U299 ( .A(n457), .B(n456), .ZN(SUM[10]) );
  NAND2_X1 U300 ( .A1(n448), .A2(n452), .ZN(n457) );
  XNOR2_X1 U301 ( .A(n319), .B(n244), .ZN(SUM[2]) );
  NAND2_X1 U302 ( .A1(n324), .A2(n243), .ZN(n319) );
  XNOR2_X1 U303 ( .A(n154), .B(n112), .ZN(SUM[5]) );
  NAND2_X1 U304 ( .A1(n111), .A2(n110), .ZN(n154) );
  XNOR2_X1 U305 ( .A(n107), .B(n105), .ZN(SUM[6]) );
  NAND2_X1 U306 ( .A1(n106), .A2(n103), .ZN(n107) );
  XNOR2_X1 U307 ( .A(n391), .B(n596), .ZN(SUM[1]) );
  NAND2_X1 U308 ( .A1(n322), .A2(n321), .ZN(n391) );
  OAI21_X1 U309 ( .B1(n465), .B2(n466), .A(n246), .ZN(n427) );
  NAND2_X1 U310 ( .A1(n324), .A2(n245), .ZN(n466) );
  NOR2_X1 U311 ( .A1(n467), .A2(n468), .ZN(n465) );
  NAND2_X1 U312 ( .A1(n243), .A2(n321), .ZN(n468) );
  OAI21_X1 U313 ( .B1(n584), .B2(n583), .A(n94), .ZN(n456) );
  INV_X1 U314 ( .A(n92), .ZN(n584) );
  OAI21_X1 U315 ( .B1(n589), .B2(n592), .A(n156), .ZN(n112) );
  INV_X1 U316 ( .A(n157), .ZN(n589) );
  OAI21_X1 U317 ( .B1(n588), .B2(n587), .A(n110), .ZN(n105) );
  INV_X1 U318 ( .A(n112), .ZN(n588) );
  INV_X1 U319 ( .A(n111), .ZN(n587) );
  OAI21_X1 U320 ( .B1(n460), .B2(n461), .A(n101), .ZN(n429) );
  NAND2_X1 U321 ( .A1(n102), .A2(n103), .ZN(n461) );
  NOR2_X1 U322 ( .A1(n15), .A2(n462), .ZN(n460) );
  AND2_X1 U323 ( .A1(n110), .A2(n156), .ZN(n15) );
  NAND4_X1 U324 ( .A1(n157), .A2(n111), .A3(n106), .A4(n101), .ZN(n430) );
  AOI21_X1 U326 ( .B1(n116), .B2(n117), .A(n118), .ZN(n113) );
  NAND2_X1 U327 ( .A1(n119), .A2(n120), .ZN(n118) );
  NOR2_X1 U328 ( .A1(n569), .A2(n570), .ZN(n116) );
  OAI211_X1 U329 ( .C1(n523), .C2(n88), .A(n122), .B(n123), .ZN(n117) );
  NOR2_X1 U331 ( .A1(n594), .A2(n392), .ZN(n467) );
  INV_X1 U333 ( .A(n322), .ZN(n594) );
  NAND2_X1 U334 ( .A1(n320), .A2(n321), .ZN(n244) );
  NAND2_X1 U335 ( .A1(n322), .A2(n596), .ZN(n320) );
  NAND2_X1 U336 ( .A1(n459), .A2(n98), .ZN(n92) );
  NAND2_X1 U337 ( .A1(n96), .A2(n97), .ZN(n459) );
  INV_X1 U338 ( .A(n392), .ZN(n596) );
  NAND2_X1 U339 ( .A1(n591), .A2(n582), .ZN(n426) );
  AND3_X1 U340 ( .A1(n93), .A2(n97), .A3(n448), .ZN(n86) );
  INV_X1 U341 ( .A(n93), .ZN(n583) );
  INV_X1 U342 ( .A(n440), .ZN(n580) );
  NAND2_X1 U343 ( .A1(n111), .A2(n106), .ZN(n462) );
  INV_X1 U344 ( .A(n324), .ZN(n593) );
  INV_X1 U345 ( .A(n115), .ZN(n568) );
  NOR2_X1 U347 ( .A1(B[60]), .A2(A[60]), .ZN(n88) );
  OR2_X1 U348 ( .A1(n530), .A2(n424), .ZN(n61) );
  AOI21_X1 U349 ( .B1(n356), .B2(n357), .A(n358), .ZN(n288) );
  AND2_X1 U350 ( .A1(n362), .A2(n363), .ZN(n356) );
  NAND2_X1 U351 ( .A1(n551), .A2(n360), .ZN(n357) );
  OAI211_X1 U352 ( .C1(n387), .C2(n388), .A(n389), .B(n390), .ZN(n386) );
  AND2_X1 U353 ( .A1(n382), .A2(n381), .ZN(n385) );
  NAND2_X1 U354 ( .A1(A[16]), .A2(B[16]), .ZN(n388) );
  NAND2_X1 U355 ( .A1(B[28]), .A2(A[28]), .ZN(n294) );
  NOR2_X1 U356 ( .A1(B[33]), .A2(A[33]), .ZN(n78) );
  NAND2_X1 U357 ( .A1(B[40]), .A2(A[40]), .ZN(net494937) );
  NAND2_X1 U358 ( .A1(A[14]), .A2(B[14]), .ZN(n413) );
  AND2_X1 U359 ( .A1(n257), .A2(n256), .ZN(n14) );
  OR2_X1 U361 ( .A1(A[35]), .A2(B[35]), .ZN(n259) );
  NAND2_X1 U362 ( .A1(B[17]), .A2(A[17]), .ZN(n398) );
  NAND2_X1 U363 ( .A1(B[12]), .A2(A[12]), .ZN(n417) );
  XNOR2_X1 U364 ( .A(n403), .B(n402), .ZN(SUM[17]) );
  OAI21_X1 U365 ( .B1(A[17]), .B2(B[17]), .A(n398), .ZN(n402) );
  NAND2_X1 U366 ( .A1(n56), .A2(n401), .ZN(n403) );
  NAND2_X1 U367 ( .A1(n52), .A2(n380), .ZN(n56) );
  OAI21_X1 U368 ( .B1(n412), .B2(n80), .A(n413), .ZN(n409) );
  AND2_X1 U369 ( .A1(n416), .A2(n417), .ZN(n80) );
  NAND2_X1 U370 ( .A1(n414), .A2(n415), .ZN(n412) );
  OR2_X1 U371 ( .A1(B[14]), .A2(A[14]), .ZN(n414) );
  NAND2_X1 U372 ( .A1(B[45]), .A2(A[45]), .ZN(net494903) );
  NAND2_X1 U373 ( .A1(A[35]), .A2(B[35]), .ZN(n262) );
  NAND2_X1 U374 ( .A1(B[22]), .A2(A[22]), .ZN(n362) );
  NAND2_X1 U375 ( .A1(B[36]), .A2(A[36]), .ZN(n236) );
  OR2_X1 U376 ( .A1(B[16]), .A2(A[16]), .ZN(n380) );
  NAND2_X1 U377 ( .A1(B[44]), .A2(A[44]), .ZN(net494902) );
  NAND2_X1 U378 ( .A1(A[10]), .A2(B[10]), .ZN(n452) );
  NAND2_X1 U379 ( .A1(A[19]), .A2(B[19]), .ZN(n286) );
  NAND2_X1 U381 ( .A1(B[34]), .A2(A[34]), .ZN(n266) );
  NAND2_X1 U382 ( .A1(B[60]), .A2(A[60]), .ZN(n123) );
  NAND2_X1 U383 ( .A1(B[57]), .A2(A[57]), .ZN(n146) );
  NOR2_X1 U384 ( .A1(A[17]), .A2(B[17]), .ZN(n387) );
  NAND2_X1 U385 ( .A1(B[62]), .A2(A[62]), .ZN(n120) );
  NAND2_X1 U386 ( .A1(B[61]), .A2(A[61]), .ZN(n122) );
  NAND2_X1 U387 ( .A1(B[18]), .A2(A[18]), .ZN(n389) );
  NAND2_X1 U388 ( .A1(B[58]), .A2(A[58]), .ZN(n147) );
  NAND2_X1 U389 ( .A1(B[21]), .A2(A[21]), .ZN(n363) );
  NAND2_X1 U390 ( .A1(B[46]), .A2(A[46]), .ZN(net494904) );
  NAND2_X1 U391 ( .A1(B[56]), .A2(A[56]), .ZN(n145) );
  NAND2_X1 U392 ( .A1(B[16]), .A2(A[16]), .ZN(n401) );
  NAND2_X1 U393 ( .A1(B[32]), .A2(A[32]), .ZN(n264) );
  NAND2_X1 U394 ( .A1(B[13]), .A2(A[13]), .ZN(n416) );
  NAND2_X1 U395 ( .A1(B[42]), .A2(A[42]), .ZN(net494931) );
  NAND2_X1 U396 ( .A1(B[48]), .A2(A[48]), .ZN(n208) );
  NAND2_X1 U397 ( .A1(B[50]), .A2(A[50]), .ZN(n209) );
  OR2_X1 U398 ( .A1(B[10]), .A2(A[10]), .ZN(n448) );
  NAND2_X1 U399 ( .A1(B[52]), .A2(A[52]), .ZN(n177) );
  NAND2_X1 U400 ( .A1(B[54]), .A2(A[54]), .ZN(n179) );
  NAND2_X1 U401 ( .A1(B[30]), .A2(A[30]), .ZN(n296) );
  NAND2_X1 U402 ( .A1(B[29]), .A2(A[29]), .ZN(n295) );
  NAND2_X1 U403 ( .A1(B[24]), .A2(A[24]), .ZN(n353) );
  NAND2_X1 U404 ( .A1(B[33]), .A2(A[33]), .ZN(n265) );
  NAND2_X1 U405 ( .A1(B[17]), .A2(A[17]), .ZN(n390) );
  NAND2_X1 U406 ( .A1(B[20]), .A2(A[20]), .ZN(n361) );
  NAND2_X1 U407 ( .A1(B[49]), .A2(A[49]), .ZN(n210) );
  NAND2_X1 U408 ( .A1(B[63]), .A2(A[63]), .ZN(n119) );
  INV_X1 U409 ( .A(B[11]), .ZN(n591) );
  OR2_X1 U410 ( .A1(B[17]), .A2(A[17]), .ZN(n399) );
  OR2_X1 U411 ( .A1(A[14]), .A2(B[14]), .ZN(n424) );
  OR2_X1 U412 ( .A1(A[35]), .A2(B[35]), .ZN(n18) );
  OR2_X1 U413 ( .A1(B[63]), .A2(A[63]), .ZN(n115) );
  NAND2_X1 U414 ( .A1(n340), .A2(n59), .ZN(n278) );
  NOR2_X1 U415 ( .A1(n85), .A2(n341), .ZN(n340) );
  OR2_X1 U416 ( .A1(n339), .A2(n540), .ZN(n59) );
  INV_X1 U417 ( .A(B[27]), .ZN(n590) );
  OR2_X1 U418 ( .A1(B[61]), .A2(A[61]), .ZN(n133) );
  OR2_X1 U419 ( .A1(B[62]), .A2(A[62]), .ZN(n129) );
  OR2_X1 U420 ( .A1(B[57]), .A2(A[57]), .ZN(n152) );
  OR2_X1 U421 ( .A1(B[56]), .A2(A[56]), .ZN(n151) );
  OR2_X1 U422 ( .A1(B[47]), .A2(A[47]), .ZN(net494895) );
  AND2_X1 U423 ( .A1(B[55]), .A2(A[55]), .ZN(n89) );
  OR2_X1 U424 ( .A1(A[33]), .A2(B[33]), .ZN(n257) );
  OR2_X1 U425 ( .A1(B[59]), .A2(A[59]), .ZN(n153) );
  INV_X1 U426 ( .A(n37), .ZN(n534) );
  OAI21_X1 U427 ( .B1(B[21]), .B2(A[21]), .A(n365), .ZN(n37) );
  NAND2_X1 U428 ( .A1(n448), .A2(n456), .ZN(n455) );
  OR2_X1 U429 ( .A1(B[6]), .A2(A[6]), .ZN(n106) );
  OR2_X1 U430 ( .A1(B[5]), .A2(A[5]), .ZN(n111) );
  OR2_X1 U431 ( .A1(B[7]), .A2(A[7]), .ZN(n101) );
  OR2_X1 U432 ( .A1(B[1]), .A2(A[1]), .ZN(n322) );
  OR2_X1 U433 ( .A1(B[2]), .A2(A[2]), .ZN(n324) );
  OR2_X1 U434 ( .A1(B[4]), .A2(A[4]), .ZN(n157) );
  OR2_X1 U435 ( .A1(B[8]), .A2(A[8]), .ZN(n97) );
  OR2_X1 U436 ( .A1(B[9]), .A2(A[9]), .ZN(n93) );
  OR2_X1 U437 ( .A1(B[3]), .A2(A[3]), .ZN(n245) );
  OR2_X1 U438 ( .A1(B[0]), .A2(A[0]), .ZN(n464) );
  NAND2_X1 U439 ( .A1(B[1]), .A2(A[1]), .ZN(n321) );
  NAND2_X1 U440 ( .A1(B[8]), .A2(A[8]), .ZN(n98) );
  NAND2_X1 U441 ( .A1(B[9]), .A2(A[9]), .ZN(n94) );
  NAND2_X1 U442 ( .A1(B[6]), .A2(A[6]), .ZN(n103) );
  NAND2_X1 U443 ( .A1(B[2]), .A2(A[2]), .ZN(n243) );
  NAND2_X1 U444 ( .A1(B[0]), .A2(A[0]), .ZN(n392) );
  NAND2_X1 U445 ( .A1(B[4]), .A2(A[4]), .ZN(n156) );
  NAND2_X1 U446 ( .A1(B[5]), .A2(A[5]), .ZN(n110) );
  NAND2_X1 U447 ( .A1(B[3]), .A2(A[3]), .ZN(n246) );
  NAND2_X1 U448 ( .A1(B[7]), .A2(A[7]), .ZN(n102) );
  AOI21_X1 U449 ( .B1(n366), .B2(n365), .A(n551), .ZN(n373) );
  OAI21_X1 U450 ( .B1(n551), .B2(n366), .A(n534), .ZN(n47) );
  AOI21_X1 U451 ( .B1(n347), .B2(n303), .A(n540), .ZN(n344) );
  XNOR2_X1 U452 ( .A(n434), .B(n435), .ZN(SUM[14]) );
  NAND2_X1 U453 ( .A1(n385), .A2(n386), .ZN(n285) );
  OAI221_X1 U454 ( .B1(n405), .B2(n406), .C1(n405), .C2(n529), .A(n411), .ZN(
        n307) );
  OAI21_X1 U455 ( .B1(A[15]), .B2(B[15]), .A(n411), .ZN(n431) );
  NOR2_X1 U456 ( .A1(A[15]), .A2(B[15]), .ZN(n405) );
  OR2_X1 U457 ( .A1(A[15]), .A2(B[15]), .ZN(n408) );
  INV_X1 U458 ( .A(n182), .ZN(n564) );
  NOR2_X1 U459 ( .A1(A[26]), .A2(B[26]), .ZN(n341) );
  NAND2_X1 U460 ( .A1(B[26]), .A2(A[26]), .ZN(n348) );
  OAI21_X1 U461 ( .B1(n556), .B2(n489), .A(net494903), .ZN(net537812) );
  OR2_X1 U462 ( .A1(B[23]), .A2(A[23]), .ZN(n64) );
  NAND2_X1 U463 ( .A1(A[23]), .A2(B[23]), .ZN(n364) );
  NAND2_X1 U464 ( .A1(n485), .A2(n286), .ZN(n284) );
  AND2_X1 U465 ( .A1(n286), .A2(n285), .ZN(n377) );
  OAI211_X1 U466 ( .C1(n306), .C2(n528), .A(n286), .B(n285), .ZN(n27) );
  OR2_X1 U467 ( .A1(B[25]), .A2(A[25]), .ZN(n337) );
  NAND2_X1 U468 ( .A1(A[25]), .A2(B[25]), .ZN(n342) );
  NOR2_X1 U469 ( .A1(A[25]), .A2(B[25]), .ZN(n343) );
  XNOR2_X1 U470 ( .A(n135), .B(n134), .ZN(SUM[61]) );
  INV_X1 U471 ( .A(n134), .ZN(n522) );
  NAND2_X1 U472 ( .A1(B[41]), .A2(A[41]), .ZN(net494936) );
  OR2_X1 U473 ( .A1(B[51]), .A2(A[51]), .ZN(n205) );
  NAND2_X1 U474 ( .A1(n54), .A2(n499), .ZN(n249) );
  OAI21_X1 U475 ( .B1(n57), .B2(n558), .A(n235), .ZN(n54) );
  XNOR2_X1 U476 ( .A(n501), .B(n349), .ZN(SUM[26]) );
  OAI21_X1 U477 ( .B1(A[23]), .B2(B[23]), .A(n359), .ZN(n358) );
  AND2_X1 U478 ( .A1(n336), .A2(n337), .ZN(n84) );
  INV_X1 U479 ( .A(n337), .ZN(n544) );
  AOI21_X1 U480 ( .B1(n408), .B2(n409), .A(n487), .ZN(n407) );
  INV_X1 U481 ( .A(n409), .ZN(n529) );
  NAND2_X1 U482 ( .A1(n214), .A2(n204), .ZN(n213) );
  NOR2_X1 U483 ( .A1(B[55]), .A2(A[55]), .ZN(n518) );
  NAND2_X1 U484 ( .A1(A[31]), .A2(B[31]), .ZN(n292) );
  NAND4_X1 U485 ( .A1(n183), .A2(n184), .A3(n182), .A4(n185), .ZN(n171) );
  OR2_X1 U486 ( .A1(B[55]), .A2(A[55]), .ZN(n185) );
  XNOR2_X1 U487 ( .A(n131), .B(n130), .ZN(SUM[62]) );
  INV_X1 U488 ( .A(n130), .ZN(n521) );
  NAND2_X1 U489 ( .A1(B[53]), .A2(A[53]), .ZN(n178) );
  AOI21_X1 U490 ( .B1(n342), .B2(n353), .A(n343), .ZN(n339) );
  NAND2_X1 U491 ( .A1(n213), .A2(n209), .ZN(n212) );
  NAND2_X1 U492 ( .A1(n230), .A2(n229), .ZN(n247) );
  OAI21_X1 U493 ( .B1(n227), .B2(n228), .A(n229), .ZN(net494888) );
  OAI21_X1 U494 ( .B1(n66), .B2(n78), .A(n265), .ZN(n270) );
  NAND2_X1 U495 ( .A1(A[15]), .A2(B[15]), .ZN(n411) );
  NAND2_X1 U496 ( .A1(A[43]), .A2(B[43]), .ZN(net494930) );
  XNOR2_X1 U497 ( .A(n309), .B(n308), .ZN(SUM[31]) );
  OAI21_X1 U498 ( .B1(n139), .B2(n524), .A(n141), .ZN(n138) );
  NOR2_X1 U499 ( .A1(n574), .A2(n573), .ZN(n142) );
  NOR2_X1 U500 ( .A1(n574), .A2(n90), .ZN(n159) );
  XNOR2_X1 U501 ( .A(n8), .B(n7), .ZN(SUM[33]) );
  AOI21_X1 U502 ( .B1(n226), .B2(n256), .A(n559), .ZN(n66) );
  NAND2_X1 U503 ( .A1(B[37]), .A2(A[37]), .ZN(n235) );
  AOI21_X1 U504 ( .B1(n150), .B2(n160), .A(n572), .ZN(n158) );
  NAND4_X1 U505 ( .A1(n224), .A2(net535402), .A3(n555), .A4(n83), .ZN(
        net494878) );
  OAI21_X1 U506 ( .B1(net494949), .B2(n554), .A(net494936), .ZN(net537213) );
  NAND2_X1 U507 ( .A1(net494933), .A2(net494936), .ZN(net494954) );
  NAND2_X1 U508 ( .A1(net494936), .A2(net494937), .ZN(net494934) );
  OAI21_X1 U509 ( .B1(n310), .B2(n311), .A(n296), .ZN(n309) );
  OAI211_X1 U510 ( .C1(n306), .C2(n528), .A(n286), .B(n485), .ZN(n366) );
  XNOR2_X1 U511 ( .A(n367), .B(n368), .ZN(SUM[22]) );
  NAND2_X1 U512 ( .A1(n47), .A2(n363), .ZN(n367) );
  NAND2_X1 U513 ( .A1(n433), .A2(n63), .ZN(n60) );
  NAND2_X1 U514 ( .A1(n433), .A2(n416), .ZN(n435) );
  NAND4_X1 U515 ( .A1(n151), .A2(n152), .A3(n150), .A4(n153), .ZN(n139) );
  INV_X1 U516 ( .A(n153), .ZN(n574) );
  NAND2_X1 U517 ( .A1(net494922), .A2(net494892), .ZN(net494921) );
  AOI21_X1 U518 ( .B1(n174), .B2(n175), .A(n89), .ZN(n173) );
  NOR2_X1 U519 ( .A1(n564), .A2(n518), .ZN(n174) );
  NAND2_X1 U520 ( .A1(net494945), .A2(net494935), .ZN(net494944) );
  NAND2_X1 U521 ( .A1(n317), .A2(n294), .ZN(n313) );
  AOI21_X1 U522 ( .B1(n226), .B2(n256), .A(n559), .ZN(n8) );
  XNOR2_X1 U523 ( .A(n158), .B(n159), .ZN(SUM[59]) );
  AND2_X1 U524 ( .A1(B[59]), .A2(A[59]), .ZN(n90) );
  OAI21_X1 U525 ( .B1(n579), .B2(n206), .A(n207), .ZN(n198) );
  AND2_X1 U526 ( .A1(n204), .A2(n205), .ZN(n207) );
  XNOR2_X1 U527 ( .A(n520), .B(n164), .ZN(SUM[57]) );
  OAI21_X1 U528 ( .B1(n476), .B2(B[11]), .A(n443), .ZN(n453) );
  NAND2_X1 U529 ( .A1(n415), .A2(n436), .ZN(n433) );
  NAND2_X1 U530 ( .A1(B[11]), .A2(n476), .ZN(n443) );
  INV_X1 U531 ( .A(n476), .ZN(n582) );
  INV_X1 U532 ( .A(net538681), .ZN(n519) );
  XNOR2_X1 U533 ( .A(net538681), .B(net494958), .ZN(SUM[40]) );
  NAND2_X1 U534 ( .A1(net538681), .A2(net494938), .ZN(net494955) );
  NAND2_X1 U535 ( .A1(A[39]), .A2(B[39]), .ZN(n230) );
  INV_X1 U536 ( .A(net494883), .ZN(n555) );
  OAI21_X1 U537 ( .B1(net494882), .B2(n477), .A(n21), .ZN(net494881) );
  OAI21_X1 U538 ( .B1(n519), .B2(net494883), .A(n21), .ZN(net537811) );
  OAI21_X1 U539 ( .B1(net494883), .B2(n519), .A(net494884), .ZN(net494922) );
  XNOR2_X1 U540 ( .A(n394), .B(n393), .ZN(SUM[19]) );
  NAND2_X1 U541 ( .A1(n307), .A2(n380), .ZN(n400) );
  NOR2_X1 U542 ( .A1(n518), .A2(n89), .ZN(n187) );
  OAI21_X1 U543 ( .B1(n77), .B2(n544), .A(n481), .ZN(n347) );
  NAND2_X1 U544 ( .A1(n40), .A2(net494895), .ZN(n6) );
  AND2_X1 U545 ( .A1(net494895), .A2(net494894), .ZN(net494899) );
  INV_X1 U546 ( .A(n166), .ZN(n520) );
  XNOR2_X1 U547 ( .A(n376), .B(n473), .ZN(SUM[20]) );
  NAND2_X1 U548 ( .A1(n369), .A2(n70), .ZN(n67) );
  OAI21_X1 U549 ( .B1(n551), .B2(n27), .A(n534), .ZN(n369) );
  AND3_X1 U550 ( .A1(n273), .A2(n41), .A3(n275), .ZN(n75) );
  XNOR2_X1 U551 ( .A(n270), .B(n271), .ZN(SUM[34]) );
  NAND2_X1 U552 ( .A1(n270), .A2(n258), .ZN(n269) );
  INV_X1 U553 ( .A(net494888), .ZN(n553) );
  OAI21_X1 U554 ( .B1(n25), .B2(n554), .A(net494936), .ZN(net494945) );
  NAND2_X1 U555 ( .A1(n495), .A2(net494888), .ZN(net538681) );
  NAND2_X1 U556 ( .A1(net494959), .A2(net494888), .ZN(net494939) );
  NAND2_X1 U557 ( .A1(A[38]), .A2(B[38]), .ZN(n231) );
  NAND2_X1 U558 ( .A1(n83), .A2(n478), .ZN(net494959) );
  NAND2_X1 U560 ( .A1(n254), .A2(n236), .ZN(n252) );
  AOI21_X1 U562 ( .B1(n237), .B2(n238), .A(n552), .ZN(n57) );
  NAND2_X1 U563 ( .A1(n479), .A2(n238), .ZN(n254) );
  XNOR2_X1 U564 ( .A(n525), .B(n192), .ZN(SUM[53]) );
  OAI21_X1 U565 ( .B1(n525), .B2(n567), .A(n178), .ZN(n188) );
  OAI21_X1 U566 ( .B1(n79), .B2(n305), .A(n355), .ZN(n51) );
  OAI21_X1 U567 ( .B1(n79), .B2(n305), .A(n355), .ZN(n331) );
  XNOR2_X1 U568 ( .A(n314), .B(n315), .ZN(SUM[30]) );
  XNOR2_X1 U569 ( .A(n328), .B(n318), .ZN(SUM[28]) );
  AOI21_X1 U570 ( .B1(n318), .B2(n300), .A(n545), .ZN(n325) );
  NAND2_X1 U571 ( .A1(n318), .A2(n300), .ZN(n317) );
  NAND2_X1 U572 ( .A1(A[27]), .A2(B[27]), .ZN(n279) );
  INV_X1 U573 ( .A(A[27]), .ZN(n541) );
  OAI21_X1 U574 ( .B1(n405), .B2(n24), .A(n407), .ZN(n53) );
  NAND2_X1 U575 ( .A1(net494894), .A2(n39), .ZN(net494911) );
  INV_X1 U576 ( .A(n194), .ZN(n525) );
  NAND2_X1 U577 ( .A1(B[51]), .A2(A[51]), .ZN(n199) );
  OAI21_X1 U578 ( .B1(net494928), .B2(n10), .A(net494929), .ZN(net494884) );
  NAND2_X1 U579 ( .A1(net494930), .A2(net494931), .ZN(net494928) );
  OAI21_X1 U580 ( .B1(n489), .B2(n556), .A(net494903), .ZN(n39) );
  XNOR2_X1 U581 ( .A(n527), .B(n218), .ZN(SUM[49]) );
  NAND2_X1 U582 ( .A1(B[47]), .A2(A[47]), .ZN(n40) );
  OAI21_X1 U583 ( .B1(n171), .B2(n498), .A(n173), .ZN(n170) );
  XNOR2_X1 U584 ( .A(n186), .B(n187), .ZN(SUM[55]) );
  AOI21_X1 U585 ( .B1(n182), .B2(n188), .A(n565), .ZN(n186) );
  XNOR2_X1 U586 ( .A(n498), .B(n196), .ZN(SUM[52]) );
  OAI21_X1 U587 ( .B1(n563), .B2(n172), .A(n177), .ZN(n194) );
  OAI21_X1 U590 ( .B1(n30), .B2(n561), .A(n208), .ZN(n220) );
  AND4_X2 U591 ( .A1(net494876), .A2(n40), .A3(net494878), .A4(net494879), 
        .ZN(n30) );
  INV_X1 U592 ( .A(n220), .ZN(n527) );
endmodule


module RCA_NBIT64_11 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_11_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), 
        .SUM({Co, S}) );
endmodule


module RCA_NBIT64_10_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net496120, net496115, net496114, net496113, net496109, net496106,
         net496057, net496040, net496036, net496035, net496030, net496026,
         net496023, net496022, net496014, net496010, net496008, net496007,
         net496006, net496005, net495996, net495993, net495992, net495991,
         net495986, net495985, net495983, net495977, net495965, net495961,
         net495943, net495933, net495932, net495929, net534711, net537211,
         net537810, net537887, net538106, net538261, net538259, net538392,
         net538497, net495948, net495945, net495942, net495939, net495944,
         net495938, net495937, net535392, net495980, net496000, net496003,
         net496002, net496001, net538867, net495999, net495987, net495982,
         net495978, net495973, net495972, net495971, net495970, n1, n2, n5, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, n21, n22, n23, n24,
         n25, n26, n27, n30, n31, n32, n33, n38, n40, n42, n45, n46, n47, n49,
         n50, n52, n53, n57, n58, n60, n61, n62, n65, n66, n67, n68, n70, n71,
         n72, n73, n74, n76, n77, n78, n79, n80, n81, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n106, n107, n108, n109, n110, n112, n113, n114,
         n115, n118, n119, n120, n123, n124, n125, n126, n127, n128, n129,
         n131, n132, n133, n134, n135, n136, n137, n139, n140, n141, n143,
         n145, n146, n147, n150, n151, n152, n153, n154, n156, n157, n158,
         n159, n161, n162, n164, n165, n167, n169, n170, n172, n173, n174,
         n176, n177, n178, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n209, n210, n211, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n226, n227, n228,
         n229, n231, n232, n233, n235, n237, n239, n241, n243, n244, n245,
         n246, n247, n248, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n272, n274, n275, n276, n277, n279, n280, n281, n282, n283, n284,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n298,
         n299, n302, n303, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n317, n319, n320, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n333, n334, n335, n336, n338, n339, n340,
         n341, n342, n343, n344, n345, n348, n349, n351, n352, n353, n354,
         n355, n356, n357, n359, n360, n362, n364, n365, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n380, n381, n383, n384,
         n387, n388, n389, n390, n392, n393, n394, n396, n397, n399, n400,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n420, n421, n422, n423, n425, n426,
         n427, n428, n429, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560;

  NAND3_X1 U50 ( .A1(net495970), .A2(net495971), .A3(net495972), .ZN(n31) );
  OR2_X2 U55 ( .A1(B[28]), .A2(A[28]), .ZN(n269) );
  NAND3_X1 U72 ( .A1(n76), .A2(n282), .A3(n281), .ZN(n329) );
  NAND3_X1 U78 ( .A1(net496008), .A2(net496007), .A3(n218), .ZN(net495985) );
  OR2_X2 U112 ( .A1(B[46]), .A2(A[46]), .ZN(net495996) );
  NAND3_X1 U121 ( .A1(net496113), .A2(net496115), .A3(n13), .ZN(net496000) );
  OR2_X2 U177 ( .A1(A[39]), .A2(B[39]), .ZN(net496008) );
  OR2_X2 U371 ( .A1(B[25]), .A2(A[25]), .ZN(n310) );
  NAND3_X1 U545 ( .A1(n284), .A2(n283), .A3(n444), .ZN(n256) );
  NAND3_X1 U571 ( .A1(n373), .A2(n372), .A3(n371), .ZN(n368) );
  NAND3_X1 U581 ( .A1(n408), .A2(n409), .A3(n410), .ZN(n407) );
  NAND3_X1 U582 ( .A1(n411), .A2(n89), .A3(n412), .ZN(n408) );
  OR2_X2 U25 ( .A1(A[34]), .A2(B[34]), .ZN(net496115) );
  OR2_X2 U113 ( .A1(B[45]), .A2(A[45]), .ZN(net496002) );
  OR2_X2 U152 ( .A1(B[50]), .A2(A[50]), .ZN(net495945) );
  OR2_X2 U350 ( .A1(B[54]), .A2(A[54]), .ZN(n181) );
  OR2_X2 U401 ( .A1(B[48]), .A2(A[48]), .ZN(net495943) );
  CLKBUF_X1 U2 ( .A(n280), .Z(n433) );
  OR2_X1 U3 ( .A1(B[24]), .A2(A[24]), .ZN(n314) );
  OR2_X1 U4 ( .A1(B[32]), .A2(A[32]), .ZN(net496114) );
  OR2_X1 U5 ( .A1(B[29]), .A2(A[29]), .ZN(n287) );
  AND2_X1 U6 ( .A1(n425), .A2(n352), .ZN(SUM[0]) );
  AND3_X1 U7 ( .A1(n256), .A2(n257), .A3(n258), .ZN(net538392) );
  OR2_X1 U8 ( .A1(B[36]), .A2(A[36]), .ZN(net496005) );
  OR2_X1 U9 ( .A1(A[38]), .A2(B[38]), .ZN(net496007) );
  OR2_X1 U10 ( .A1(B[44]), .A2(A[44]), .ZN(net496001) );
  OR2_X1 U11 ( .A1(A[49]), .A2(B[49]), .ZN(net495944) );
  OR2_X1 U12 ( .A1(B[51]), .A2(A[51]), .ZN(net495942) );
  OR2_X1 U13 ( .A1(B[52]), .A2(A[52]), .ZN(n183) );
  OR2_X1 U14 ( .A1(B[56]), .A2(A[56]), .ZN(n151) );
  BUF_X1 U15 ( .A(n38), .Z(n434) );
  AND2_X1 U16 ( .A1(net535392), .A2(n478), .ZN(n435) );
  AOI21_X1 U17 ( .B1(net495932), .B2(net495933), .A(n517), .ZN(n436) );
  INV_X1 U18 ( .A(n495), .ZN(n437) );
  CLKBUF_X1 U19 ( .A(A[19]), .Z(n438) );
  OAI21_X1 U20 ( .B1(n481), .B2(n274), .A(n275), .ZN(n439) );
  NAND2_X1 U21 ( .A1(net537887), .A2(n241), .ZN(n440) );
  CLKBUF_X1 U22 ( .A(n205), .Z(n441) );
  OAI21_X1 U23 ( .B1(n334), .B2(n85), .A(n335), .ZN(n442) );
  AND4_X1 U24 ( .A1(n307), .A2(n450), .A3(n314), .A4(n310), .ZN(n443) );
  OR2_X1 U26 ( .A1(A[31]), .A2(B[31]), .ZN(n444) );
  OR2_X1 U27 ( .A1(A[31]), .A2(B[31]), .ZN(n267) );
  OR2_X1 U28 ( .A1(B[33]), .A2(A[33]), .ZN(n445) );
  OR2_X1 U29 ( .A1(B[33]), .A2(A[33]), .ZN(net496109) );
  AND2_X1 U30 ( .A1(n447), .A2(n448), .ZN(n446) );
  NAND2_X1 U31 ( .A1(n66), .A2(n345), .ZN(n447) );
  NAND2_X1 U32 ( .A1(n447), .A2(n448), .ZN(n57) );
  AND2_X1 U33 ( .A1(n76), .A2(n282), .ZN(n448) );
  AND3_X1 U34 ( .A1(net495970), .A2(net495971), .A3(net495972), .ZN(net538259)
         );
  OR2_X1 U35 ( .A1(B[43]), .A2(A[43]), .ZN(net496030) );
  CLKBUF_X1 U36 ( .A(n521), .Z(n449) );
  OR2_X1 U37 ( .A1(A[30]), .A2(B[30]), .ZN(n272) );
  AND2_X1 U38 ( .A1(n185), .A2(n181), .ZN(n173) );
  OR2_X1 U39 ( .A1(B[26]), .A2(A[26]), .ZN(n450) );
  NOR2_X1 U40 ( .A1(A[47]), .A2(B[47]), .ZN(n451) );
  OR2_X1 U41 ( .A1(A[47]), .A2(B[47]), .ZN(net496003) );
  INV_X1 U42 ( .A(n499), .ZN(n452) );
  OR2_X1 U43 ( .A1(A[37]), .A2(B[37]), .ZN(net496006) );
  OR2_X1 U44 ( .A1(n72), .A2(n73), .ZN(net496057) );
  OR2_X1 U45 ( .A1(B[55]), .A2(A[55]), .ZN(n185) );
  OR2_X1 U46 ( .A1(A[26]), .A2(B[26]), .ZN(n311) );
  OR2_X2 U47 ( .A1(A[16]), .A2(B[16]), .ZN(n341) );
  CLKBUF_X1 U48 ( .A(A[26]), .Z(n453) );
  AND2_X1 U49 ( .A1(n13), .A2(net496115), .ZN(n454) );
  OR2_X2 U51 ( .A1(A[17]), .A2(B[17]), .ZN(n342) );
  NAND3_X1 U52 ( .A1(net495999), .A2(n21), .A3(n435), .ZN(net495970) );
  XNOR2_X1 U53 ( .A(n440), .B(n455), .ZN(SUM[36]) );
  NAND2_X1 U54 ( .A1(net496005), .A2(n219), .ZN(n455) );
  XNOR2_X1 U56 ( .A(n465), .B(n456), .ZN(SUM[43]) );
  NAND2_X1 U57 ( .A1(n202), .A2(net496030), .ZN(n456) );
  OR2_X1 U58 ( .A1(A[42]), .A2(B[42]), .ZN(net496036) );
  OAI21_X1 U59 ( .B1(n501), .B2(n475), .A(n145), .ZN(n457) );
  NAND2_X1 U60 ( .A1(n454), .A2(net496113), .ZN(n8) );
  OR2_X1 U61 ( .A1(B[40]), .A2(A[40]), .ZN(net496040) );
  AND2_X1 U62 ( .A1(n77), .A2(net496008), .ZN(n458) );
  AND2_X1 U63 ( .A1(n458), .A2(n65), .ZN(n459) );
  OR2_X1 U64 ( .A1(A[41]), .A2(B[41]), .ZN(net496035) );
  AND2_X1 U65 ( .A1(net495942), .A2(net495945), .ZN(net495932) );
  OAI21_X1 U66 ( .B1(n470), .B2(net495980), .A(n437), .ZN(n460) );
  XNOR2_X1 U67 ( .A(n81), .B(n461), .ZN(SUM[26]) );
  NAND2_X1 U68 ( .A1(n450), .A2(n52), .ZN(n461) );
  XNOR2_X1 U69 ( .A(n462), .B(n463), .ZN(SUM[45]) );
  AND2_X1 U70 ( .A1(net496022), .A2(net495991), .ZN(n462) );
  AND2_X1 U71 ( .A1(net496002), .A2(net495992), .ZN(n463) );
  XOR2_X1 U73 ( .A(n464), .B(net537810), .Z(SUM[50]) );
  AND2_X1 U74 ( .A1(net495945), .A2(net495939), .ZN(n464) );
  NAND2_X1 U75 ( .A1(n209), .A2(n203), .ZN(n465) );
  NOR2_X1 U76 ( .A1(n486), .A2(n488), .ZN(n255) );
  INV_X1 U77 ( .A(n135), .ZN(n474) );
  NAND2_X1 U79 ( .A1(n365), .A2(n364), .ZN(n283) );
  NAND2_X1 U80 ( .A1(n80), .A2(n283), .ZN(n76) );
  AND2_X1 U81 ( .A1(n365), .A2(n364), .ZN(n58) );
  NAND2_X1 U82 ( .A1(net535392), .A2(net495982), .ZN(n45) );
  NAND2_X1 U83 ( .A1(net495983), .A2(n522), .ZN(net495982) );
  OAI21_X1 U84 ( .B1(n555), .B2(n380), .A(n389), .ZN(n92) );
  NAND2_X1 U85 ( .A1(n405), .A2(n387), .ZN(n403) );
  NAND2_X1 U86 ( .A1(n545), .A2(n92), .ZN(n405) );
  INV_X1 U87 ( .A(n390), .ZN(n545) );
  AOI21_X1 U88 ( .B1(n109), .B2(n110), .A(n507), .ZN(SUM[64]) );
  INV_X1 U89 ( .A(n392), .ZN(n555) );
  NAND2_X1 U90 ( .A1(n549), .A2(n392), .ZN(n388) );
  INV_X1 U91 ( .A(n380), .ZN(n549) );
  INV_X1 U92 ( .A(n143), .ZN(n504) );
  XNOR2_X1 U93 ( .A(n251), .B(n252), .ZN(SUM[34]) );
  NOR2_X1 U94 ( .A1(n524), .A2(n523), .ZN(n252) );
  AOI21_X1 U95 ( .B1(n254), .B2(n445), .A(n519), .ZN(n251) );
  INV_X1 U96 ( .A(net496115), .ZN(n523) );
  NAND2_X1 U97 ( .A1(n326), .A2(n325), .ZN(n333) );
  NAND2_X1 U98 ( .A1(n269), .A2(n264), .ZN(n303) );
  NAND2_X1 U99 ( .A1(net496040), .A2(n206), .ZN(n215) );
  NAND2_X1 U100 ( .A1(net496036), .A2(n203), .ZN(n211) );
  NAND2_X1 U101 ( .A1(net496001), .A2(net495991), .ZN(net496026) );
  NAND2_X1 U102 ( .A1(n131), .A2(n119), .ZN(n133) );
  NAND2_X1 U103 ( .A1(n118), .A2(n124), .ZN(n129) );
  NAND2_X1 U104 ( .A1(n266), .A2(n272), .ZN(n291) );
  NAND2_X1 U105 ( .A1(n183), .A2(n176), .ZN(n195) );
  NAND2_X1 U106 ( .A1(net495944), .A2(net495938), .ZN(net495961) );
  NAND2_X1 U107 ( .A1(n314), .A2(n313), .ZN(n320) );
  NAND2_X1 U108 ( .A1(n287), .A2(n265), .ZN(n299) );
  INV_X1 U109 ( .A(n269), .ZN(n533) );
  NAND2_X1 U110 ( .A1(n373), .A2(n369), .ZN(n397) );
  XOR2_X1 U111 ( .A(n231), .B(n466), .Z(SUM[39]) );
  AND2_X1 U114 ( .A1(net496008), .A2(net495986), .ZN(n466) );
  AOI21_X1 U115 ( .B1(net496014), .B2(net495996), .A(n492), .ZN(n198) );
  INV_X1 U116 ( .A(net495993), .ZN(n492) );
  NAND2_X1 U117 ( .A1(n282), .A2(n344), .ZN(n353) );
  INV_X1 U118 ( .A(n343), .ZN(n485) );
  NAND2_X1 U119 ( .A1(net495996), .A2(net495993), .ZN(n199) );
  XNOR2_X1 U120 ( .A(n330), .B(n79), .ZN(SUM[23]) );
  NOR2_X1 U122 ( .A1(n27), .A2(n531), .ZN(n79) );
  INV_X1 U123 ( .A(n327), .ZN(n531) );
  INV_X1 U124 ( .A(n49), .ZN(n517) );
  INV_X1 U125 ( .A(n287), .ZN(n534) );
  INV_X1 U126 ( .A(n264), .ZN(n532) );
  INV_X1 U127 ( .A(n341), .ZN(n484) );
  AND2_X1 U128 ( .A1(n310), .A2(n312), .ZN(n84) );
  AND2_X1 U129 ( .A1(n447), .A2(n282), .ZN(n14) );
  INV_X1 U130 ( .A(n27), .ZN(n530) );
  OAI21_X1 U131 ( .B1(n488), .B2(net538392), .A(net496106), .ZN(n254) );
  INV_X1 U132 ( .A(n362), .ZN(n483) );
  OAI211_X1 U133 ( .C1(n520), .C2(net496106), .A(n245), .B(n244), .ZN(n243) );
  INV_X1 U134 ( .A(net496109), .ZN(n520) );
  XNOR2_X1 U135 ( .A(n289), .B(n288), .ZN(SUM[31]) );
  NAND2_X1 U136 ( .A1(n262), .A2(n444), .ZN(n288) );
  NAND2_X1 U137 ( .A1(n290), .A2(n266), .ZN(n289) );
  XNOR2_X1 U138 ( .A(n356), .B(n355), .ZN(SUM[18]) );
  NAND2_X1 U139 ( .A1(n343), .A2(n349), .ZN(n356) );
  NOR2_X1 U140 ( .A1(n367), .A2(n539), .ZN(n365) );
  INV_X1 U141 ( .A(n376), .ZN(n539) );
  AOI22_X1 U142 ( .A1(n369), .A2(n368), .B1(n538), .B2(n559), .ZN(n367) );
  XNOR2_X1 U143 ( .A(n340), .B(n57), .ZN(SUM[20]) );
  NAND2_X1 U144 ( .A1(n339), .A2(n328), .ZN(n340) );
  XNOR2_X1 U145 ( .A(n60), .B(n233), .ZN(SUM[38]) );
  NOR2_X1 U146 ( .A1(n490), .A2(n491), .ZN(n233) );
  INV_X1 U147 ( .A(n220), .ZN(n490) );
  XOR2_X1 U148 ( .A(n58), .B(n467), .Z(SUM[16]) );
  NAND2_X1 U149 ( .A1(n341), .A2(n362), .ZN(n467) );
  XOR2_X1 U150 ( .A(n468), .B(n239), .Z(SUM[37]) );
  AND2_X1 U151 ( .A1(net496006), .A2(n221), .ZN(n468) );
  XNOR2_X1 U153 ( .A(n125), .B(n126), .ZN(SUM[63]) );
  NAND2_X1 U154 ( .A1(n123), .A2(n112), .ZN(n125) );
  XNOR2_X1 U155 ( .A(n254), .B(n253), .ZN(SUM[33]) );
  NAND2_X1 U156 ( .A1(n445), .A2(n244), .ZN(n253) );
  XNOR2_X1 U157 ( .A(n7), .B(n336), .ZN(SUM[21]) );
  NOR2_X1 U158 ( .A1(n85), .A2(n528), .ZN(n336) );
  INV_X1 U159 ( .A(n335), .ZN(n528) );
  INV_X1 U160 ( .A(net496000), .ZN(n489) );
  OAI211_X1 U161 ( .C1(n511), .C2(n176), .A(n177), .B(n178), .ZN(n174) );
  OAI21_X1 U162 ( .B1(n477), .B2(n518), .A(net495939), .ZN(n50) );
  AOI21_X1 U163 ( .B1(net495987), .B2(n46), .A(net534711), .ZN(net495971) );
  OAI211_X1 U164 ( .C1(n494), .C2(net495991), .A(net495992), .B(net495993), 
        .ZN(n46) );
  INV_X1 U165 ( .A(net495996), .ZN(n493) );
  OAI21_X1 U166 ( .B1(n473), .B2(n509), .A(n119), .ZN(n128) );
  OAI21_X1 U167 ( .B1(n334), .B2(n85), .A(n335), .ZN(n53) );
  INV_X1 U168 ( .A(n178), .ZN(n513) );
  INV_X1 U169 ( .A(n177), .ZN(n510) );
  XNOR2_X1 U170 ( .A(n136), .B(n135), .ZN(SUM[60]) );
  NAND2_X1 U171 ( .A1(n134), .A2(n120), .ZN(n136) );
  XNOR2_X1 U172 ( .A(n246), .B(net496120), .ZN(SUM[35]) );
  NAND2_X1 U173 ( .A1(n445), .A2(net496115), .ZN(n247) );
  OAI21_X1 U174 ( .B1(n201), .B2(n200), .A(net496030), .ZN(net495977) );
  AND3_X1 U175 ( .A1(net496035), .A2(net496036), .A3(n204), .ZN(n200) );
  OAI21_X1 U176 ( .B1(net495973), .B2(n495), .A(net538867), .ZN(net495972) );
  AOI21_X1 U178 ( .B1(net495978), .B2(n45), .A(net495980), .ZN(net495973) );
  OR2_X1 U179 ( .A1(net496000), .A2(n23), .ZN(net537887) );
  OAI21_X1 U180 ( .B1(net538106), .B2(n494), .A(net495992), .ZN(net496014) );
  AOI21_X1 U181 ( .B1(net496115), .B2(n519), .A(n524), .ZN(n248) );
  NAND4_X1 U182 ( .A1(n268), .A2(n269), .A3(n444), .A4(n270), .ZN(n257) );
  OAI21_X1 U183 ( .B1(n479), .B2(n274), .A(n19), .ZN(n268) );
  AND2_X1 U184 ( .A1(n287), .A2(n272), .ZN(n270) );
  INV_X1 U185 ( .A(n276), .ZN(n479) );
  OAI211_X1 U186 ( .C1(n502), .C2(n145), .A(n146), .B(n147), .ZN(n141) );
  NOR2_X1 U187 ( .A1(n309), .A2(n78), .ZN(n305) );
  AND2_X1 U188 ( .A1(n312), .A2(n313), .ZN(n78) );
  NAND2_X1 U189 ( .A1(n311), .A2(n310), .ZN(n309) );
  AND4_X1 U190 ( .A1(n287), .A2(n272), .A3(n15), .A4(n26), .ZN(n284) );
  AND2_X1 U191 ( .A1(n526), .A2(n269), .ZN(n15) );
  AND2_X1 U192 ( .A1(n443), .A2(n80), .ZN(n26) );
  OAI21_X1 U193 ( .B1(n544), .B2(n543), .A(n375), .ZN(n399) );
  INV_X1 U194 ( .A(n403), .ZN(n544) );
  NAND2_X1 U195 ( .A1(n216), .A2(net496005), .ZN(n237) );
  OAI211_X1 U196 ( .C1(n499), .C2(n219), .A(n220), .B(n221), .ZN(n218) );
  OAI21_X1 U197 ( .B1(n317), .B2(n537), .A(n312), .ZN(n315) );
  NOR2_X1 U198 ( .A1(n500), .A2(n501), .ZN(n167) );
  INV_X1 U199 ( .A(n145), .ZN(n500) );
  INV_X1 U200 ( .A(net496002), .ZN(n494) );
  AND3_X1 U201 ( .A1(n344), .A2(n5), .A3(n343), .ZN(n80) );
  INV_X1 U202 ( .A(A[15]), .ZN(n538) );
  INV_X1 U203 ( .A(n40), .ZN(n522) );
  AND3_X1 U204 ( .A1(net496008), .A2(n65), .A3(n77), .ZN(n73) );
  AND2_X1 U205 ( .A1(net496007), .A2(n217), .ZN(n77) );
  OAI21_X1 U206 ( .B1(n71), .B2(n496), .A(n206), .ZN(n213) );
  NOR2_X1 U207 ( .A1(n459), .A2(n72), .ZN(n71) );
  INV_X1 U208 ( .A(n245), .ZN(n524) );
  INV_X1 U209 ( .A(n244), .ZN(n519) );
  INV_X1 U210 ( .A(n373), .ZN(n540) );
  INV_X1 U211 ( .A(n131), .ZN(n509) );
  INV_X1 U212 ( .A(n184), .ZN(n511) );
  NAND2_X1 U213 ( .A1(n308), .A2(n52), .ZN(n306) );
  INV_X1 U214 ( .A(net496114), .ZN(n488) );
  AND3_X1 U215 ( .A1(n256), .A2(n2), .A3(n257), .ZN(n23) );
  AND2_X1 U216 ( .A1(net496022), .A2(net495991), .ZN(net538106) );
  INV_X1 U217 ( .A(n310), .ZN(n537) );
  INV_X1 U218 ( .A(net496106), .ZN(n486) );
  INV_X1 U219 ( .A(net495944), .ZN(n516) );
  AND3_X1 U220 ( .A1(net496036), .A2(net496035), .A3(net496040), .ZN(n47) );
  INV_X1 U221 ( .A(net496040), .ZN(n496) );
  INV_X1 U222 ( .A(net495945), .ZN(n518) );
  INV_X1 U223 ( .A(net496007), .ZN(n491) );
  AND2_X1 U224 ( .A1(n194), .A2(n176), .ZN(n191) );
  INV_X1 U225 ( .A(n134), .ZN(n506) );
  INV_X1 U226 ( .A(n151), .ZN(n501) );
  NAND2_X1 U227 ( .A1(n237), .A2(n219), .ZN(n235) );
  AND2_X1 U228 ( .A1(net496109), .A2(net496114), .ZN(n13) );
  NAND2_X1 U229 ( .A1(n374), .A2(n375), .ZN(n372) );
  INV_X1 U230 ( .A(n313), .ZN(n536) );
  INV_X1 U231 ( .A(n221), .ZN(n498) );
  INV_X1 U232 ( .A(n262), .ZN(n535) );
  INV_X1 U233 ( .A(net496035), .ZN(n497) );
  INV_X1 U234 ( .A(n325), .ZN(n527) );
  AND2_X1 U235 ( .A1(net496002), .A2(net496001), .ZN(n10) );
  XNOR2_X1 U236 ( .A(n400), .B(n399), .ZN(SUM[13]) );
  NAND2_X1 U237 ( .A1(n371), .A2(n374), .ZN(n400) );
  XNOR2_X1 U238 ( .A(n95), .B(n96), .ZN(SUM[7]) );
  NAND2_X1 U239 ( .A1(n99), .A2(n100), .ZN(n95) );
  NAND2_X1 U240 ( .A1(n97), .A2(n98), .ZN(n96) );
  NAND2_X1 U241 ( .A1(n101), .A2(n102), .ZN(n100) );
  XNOR2_X1 U242 ( .A(n413), .B(n414), .ZN(SUM[11]) );
  NAND2_X1 U243 ( .A1(n409), .A2(n415), .ZN(n414) );
  NAND2_X1 U244 ( .A1(n410), .A2(n406), .ZN(n413) );
  NAND2_X1 U245 ( .A1(n412), .A2(n416), .ZN(n415) );
  XNOR2_X1 U246 ( .A(n404), .B(n403), .ZN(SUM[12]) );
  NAND2_X1 U247 ( .A1(n402), .A2(n375), .ZN(n404) );
  XNOR2_X1 U248 ( .A(n91), .B(n92), .ZN(SUM[8]) );
  NAND2_X1 U249 ( .A1(n93), .A2(n94), .ZN(n91) );
  XNOR2_X1 U250 ( .A(n293), .B(n227), .ZN(SUM[2]) );
  NAND2_X1 U251 ( .A1(n298), .A2(n226), .ZN(n293) );
  XNOR2_X1 U252 ( .A(n87), .B(n88), .ZN(SUM[9]) );
  NAND2_X1 U253 ( .A1(n89), .A2(n90), .ZN(n87) );
  XNOR2_X1 U254 ( .A(n154), .B(n108), .ZN(SUM[5]) );
  NAND2_X1 U255 ( .A1(n107), .A2(n106), .ZN(n154) );
  XNOR2_X1 U256 ( .A(n103), .B(n101), .ZN(SUM[6]) );
  NAND2_X1 U257 ( .A1(n102), .A2(n99), .ZN(n103) );
  XNOR2_X1 U258 ( .A(n417), .B(n416), .ZN(SUM[10]) );
  NAND2_X1 U259 ( .A1(n412), .A2(n409), .ZN(n417) );
  XNOR2_X1 U260 ( .A(n351), .B(n560), .ZN(SUM[1]) );
  NAND2_X1 U261 ( .A1(n296), .A2(n295), .ZN(n351) );
  XNOR2_X1 U262 ( .A(n197), .B(n392), .ZN(SUM[4]) );
  NAND2_X1 U263 ( .A1(n157), .A2(n156), .ZN(n197) );
  XNOR2_X1 U264 ( .A(n222), .B(n223), .ZN(SUM[3]) );
  OAI21_X1 U265 ( .B1(n558), .B2(n556), .A(n226), .ZN(n223) );
  NAND2_X1 U266 ( .A1(n228), .A2(n229), .ZN(n222) );
  INV_X1 U267 ( .A(n227), .ZN(n558) );
  OAI21_X1 U268 ( .B1(n426), .B2(n427), .A(n229), .ZN(n392) );
  NAND2_X1 U269 ( .A1(n298), .A2(n228), .ZN(n427) );
  NOR2_X1 U270 ( .A1(n428), .A2(n429), .ZN(n426) );
  NAND2_X1 U271 ( .A1(n226), .A2(n295), .ZN(n429) );
  OAI21_X1 U272 ( .B1(n548), .B2(n547), .A(n90), .ZN(n416) );
  INV_X1 U273 ( .A(n88), .ZN(n548) );
  INV_X1 U274 ( .A(n89), .ZN(n547) );
  OAI21_X1 U275 ( .B1(n552), .B2(n555), .A(n156), .ZN(n108) );
  INV_X1 U276 ( .A(n157), .ZN(n552) );
  OAI21_X1 U277 ( .B1(n551), .B2(n550), .A(n106), .ZN(n101) );
  INV_X1 U278 ( .A(n108), .ZN(n551) );
  INV_X1 U279 ( .A(n107), .ZN(n550) );
  NOR3_X1 U280 ( .A1(n540), .A2(n543), .A3(n1), .ZN(n384) );
  OAI21_X1 U281 ( .B1(n421), .B2(n422), .A(n97), .ZN(n389) );
  NAND2_X1 U282 ( .A1(n98), .A2(n99), .ZN(n422) );
  NOR2_X1 U283 ( .A1(n16), .A2(n423), .ZN(n421) );
  AND2_X1 U284 ( .A1(n106), .A2(n156), .ZN(n16) );
  OAI211_X1 U285 ( .C1(n381), .C2(n546), .A(n370), .B(n384), .ZN(n364) );
  INV_X1 U286 ( .A(n387), .ZN(n546) );
  NAND2_X1 U287 ( .A1(n559), .A2(n538), .ZN(n370) );
  AOI21_X1 U288 ( .B1(n388), .B2(n389), .A(n390), .ZN(n381) );
  NAND4_X1 U289 ( .A1(n157), .A2(n107), .A3(n102), .A4(n97), .ZN(n380) );
  NAND4_X1 U290 ( .A1(n89), .A2(n93), .A3(n412), .A4(n406), .ZN(n390) );
  OAI21_X1 U291 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  NAND2_X1 U292 ( .A1(n119), .A2(n120), .ZN(n114) );
  NOR2_X1 U293 ( .A1(n474), .A2(n506), .ZN(n113) );
  NOR2_X1 U294 ( .A1(n508), .A2(n509), .ZN(n115) );
  NOR2_X1 U295 ( .A1(n557), .A2(n352), .ZN(n428) );
  INV_X1 U296 ( .A(n296), .ZN(n557) );
  NAND2_X1 U297 ( .A1(n420), .A2(n94), .ZN(n88) );
  NAND2_X1 U298 ( .A1(n92), .A2(n93), .ZN(n420) );
  NAND2_X1 U299 ( .A1(n294), .A2(n295), .ZN(n227) );
  NAND2_X1 U300 ( .A1(n296), .A2(n560), .ZN(n294) );
  NAND2_X1 U301 ( .A1(n406), .A2(n407), .ZN(n387) );
  NAND2_X1 U302 ( .A1(n90), .A2(n94), .ZN(n411) );
  INV_X1 U303 ( .A(n352), .ZN(n560) );
  INV_X1 U304 ( .A(n402), .ZN(n543) );
  NAND2_X1 U305 ( .A1(n107), .A2(n102), .ZN(n423) );
  AND2_X1 U306 ( .A1(n123), .A2(n124), .ZN(n109) );
  INV_X1 U307 ( .A(n298), .ZN(n556) );
  INV_X1 U308 ( .A(n118), .ZN(n508) );
  INV_X1 U309 ( .A(n112), .ZN(n507) );
  NAND2_X1 U310 ( .A1(A[20]), .A2(B[20]), .ZN(n324) );
  NOR2_X1 U311 ( .A1(A[21]), .A2(B[21]), .ZN(n323) );
  AND2_X1 U312 ( .A1(n308), .A2(n74), .ZN(n33) );
  NAND2_X1 U313 ( .A1(n383), .A2(n376), .ZN(n393) );
  OAI21_X1 U314 ( .B1(n541), .B2(n540), .A(n369), .ZN(n394) );
  OR2_X1 U315 ( .A1(B[15]), .A2(A[15]), .ZN(n383) );
  NOR2_X1 U316 ( .A1(B[21]), .A2(A[21]), .ZN(n85) );
  NAND4_X1 U317 ( .A1(n307), .A2(n450), .A3(n314), .A4(n310), .ZN(n274) );
  OR2_X1 U318 ( .A1(B[27]), .A2(A[27]), .ZN(n307) );
  AOI22_X1 U319 ( .A1(n554), .A2(n525), .B1(n529), .B2(n553), .ZN(n83) );
  INV_X1 U320 ( .A(B[23]), .ZN(n553) );
  INV_X1 U321 ( .A(A[23]), .ZN(n529) );
  NAND4_X1 U322 ( .A1(n327), .A2(n11), .A3(n326), .A4(n328), .ZN(n277) );
  OR2_X1 U323 ( .A1(A[21]), .A2(B[21]), .ZN(n11) );
  OAI211_X1 U324 ( .C1(n263), .C2(n264), .A(n265), .B(n266), .ZN(n260) );
  NOR2_X1 U325 ( .A1(A[29]), .A2(B[29]), .ZN(n263) );
  NOR2_X1 U326 ( .A1(A[13]), .A2(B[13]), .ZN(n1) );
  NAND2_X1 U327 ( .A1(B[36]), .A2(A[36]), .ZN(n219) );
  NAND2_X1 U328 ( .A1(B[28]), .A2(A[28]), .ZN(n264) );
  NAND2_X1 U329 ( .A1(B[44]), .A2(A[44]), .ZN(net495991) );
  NAND2_X1 U330 ( .A1(B[40]), .A2(A[40]), .ZN(n206) );
  NAND2_X1 U331 ( .A1(B[45]), .A2(A[45]), .ZN(net495992) );
  NAND2_X1 U332 ( .A1(B[21]), .A2(A[21]), .ZN(n335) );
  NAND2_X1 U333 ( .A1(B[33]), .A2(A[33]), .ZN(n244) );
  NAND2_X1 U334 ( .A1(B[12]), .A2(A[12]), .ZN(n375) );
  NAND2_X1 U335 ( .A1(B[46]), .A2(A[46]), .ZN(net495993) );
  NAND2_X1 U336 ( .A1(B[61]), .A2(A[61]), .ZN(n119) );
  NAND2_X1 U337 ( .A1(B[32]), .A2(A[32]), .ZN(net496106) );
  NAND2_X1 U338 ( .A1(B[29]), .A2(A[29]), .ZN(n265) );
  NAND2_X1 U339 ( .A1(A[34]), .A2(B[34]), .ZN(n245) );
  NAND2_X1 U340 ( .A1(B[13]), .A2(A[13]), .ZN(n374) );
  NAND2_X1 U341 ( .A1(B[25]), .A2(A[25]), .ZN(n312) );
  NAND2_X1 U342 ( .A1(B[54]), .A2(A[54]), .ZN(n178) );
  NAND2_X1 U343 ( .A1(B[24]), .A2(A[24]), .ZN(n313) );
  NAND2_X1 U344 ( .A1(A[42]), .A2(B[42]), .ZN(n203) );
  NAND2_X1 U345 ( .A1(B[52]), .A2(A[52]), .ZN(n176) );
  NAND2_X1 U346 ( .A1(A[15]), .A2(B[15]), .ZN(n376) );
  NAND2_X1 U347 ( .A1(B[50]), .A2(A[50]), .ZN(net495939) );
  NAND2_X1 U348 ( .A1(B[38]), .A2(A[38]), .ZN(n220) );
  OR2_X1 U349 ( .A1(B[18]), .A2(A[18]), .ZN(n343) );
  NAND2_X1 U351 ( .A1(B[56]), .A2(A[56]), .ZN(n145) );
  NAND2_X1 U352 ( .A1(A[16]), .A2(B[16]), .ZN(n362) );
  NAND2_X1 U353 ( .A1(B[37]), .A2(A[37]), .ZN(n221) );
  OR2_X1 U354 ( .A1(B[20]), .A2(A[20]), .ZN(n328) );
  NAND2_X1 U355 ( .A1(B[41]), .A2(A[41]), .ZN(n205) );
  AND2_X1 U356 ( .A1(A[23]), .A2(B[23]), .ZN(n27) );
  NAND2_X1 U357 ( .A1(B[20]), .A2(A[20]), .ZN(n339) );
  NAND2_X1 U358 ( .A1(B[62]), .A2(A[62]), .ZN(n124) );
  NAND2_X1 U359 ( .A1(B[18]), .A2(A[18]), .ZN(n349) );
  NAND2_X1 U360 ( .A1(B[58]), .A2(A[58]), .ZN(n147) );
  INV_X1 U361 ( .A(B[15]), .ZN(n559) );
  NAND2_X1 U362 ( .A1(A[27]), .A2(B[27]), .ZN(n308) );
  OR2_X1 U363 ( .A1(B[62]), .A2(A[62]), .ZN(n118) );
  NAND2_X1 U364 ( .A1(A[31]), .A2(B[31]), .ZN(n262) );
  OR2_X1 U365 ( .A1(A[14]), .A2(B[14]), .ZN(n373) );
  NAND2_X1 U366 ( .A1(n66), .A2(n345), .ZN(n281) );
  AND2_X1 U367 ( .A1(n343), .A2(n344), .ZN(n66) );
  OR2_X1 U368 ( .A1(A[19]), .A2(B[19]), .ZN(n344) );
  INV_X1 U369 ( .A(B[22]), .ZN(n554) );
  OR2_X1 U370 ( .A1(B[63]), .A2(A[63]), .ZN(n112) );
  OR2_X1 U372 ( .A1(B[61]), .A2(A[61]), .ZN(n131) );
  OR2_X1 U373 ( .A1(A[23]), .A2(B[23]), .ZN(n327) );
  OR2_X1 U374 ( .A1(B[60]), .A2(A[60]), .ZN(n134) );
  OR2_X1 U375 ( .A1(A[27]), .A2(B[27]), .ZN(n74) );
  OR2_X1 U376 ( .A1(B[59]), .A2(A[59]), .ZN(n150) );
  OR2_X1 U377 ( .A1(B[58]), .A2(A[58]), .ZN(n153) );
  OR2_X1 U378 ( .A1(A[35]), .A2(B[35]), .ZN(net496113) );
  OR2_X1 U379 ( .A1(B[53]), .A2(A[53]), .ZN(n184) );
  OR2_X1 U380 ( .A1(A[13]), .A2(B[13]), .ZN(n371) );
  AND2_X1 U381 ( .A1(n267), .A2(n32), .ZN(n259) );
  OR2_X1 U382 ( .A1(B[6]), .A2(A[6]), .ZN(n102) );
  OR2_X1 U383 ( .A1(B[5]), .A2(A[5]), .ZN(n107) );
  OR2_X1 U384 ( .A1(B[10]), .A2(A[10]), .ZN(n412) );
  OR2_X1 U385 ( .A1(B[9]), .A2(A[9]), .ZN(n89) );
  OR2_X1 U386 ( .A1(B[11]), .A2(A[11]), .ZN(n406) );
  OR2_X1 U387 ( .A1(B[7]), .A2(A[7]), .ZN(n97) );
  OR2_X1 U388 ( .A1(B[8]), .A2(A[8]), .ZN(n93) );
  OR2_X1 U389 ( .A1(B[1]), .A2(A[1]), .ZN(n296) );
  OR2_X1 U390 ( .A1(B[2]), .A2(A[2]), .ZN(n298) );
  OR2_X1 U391 ( .A1(B[4]), .A2(A[4]), .ZN(n157) );
  OR2_X1 U392 ( .A1(B[3]), .A2(A[3]), .ZN(n228) );
  OR2_X1 U393 ( .A1(B[12]), .A2(A[12]), .ZN(n402) );
  OR2_X1 U394 ( .A1(B[0]), .A2(A[0]), .ZN(n425) );
  NAND2_X1 U395 ( .A1(B[1]), .A2(A[1]), .ZN(n295) );
  NAND2_X1 U396 ( .A1(B[8]), .A2(A[8]), .ZN(n94) );
  NAND2_X1 U397 ( .A1(B[6]), .A2(A[6]), .ZN(n99) );
  NAND2_X1 U398 ( .A1(B[9]), .A2(A[9]), .ZN(n90) );
  NAND2_X1 U399 ( .A1(B[2]), .A2(A[2]), .ZN(n226) );
  NAND2_X1 U400 ( .A1(B[0]), .A2(A[0]), .ZN(n352) );
  NAND2_X1 U402 ( .A1(B[4]), .A2(A[4]), .ZN(n156) );
  NAND2_X1 U403 ( .A1(B[5]), .A2(A[5]), .ZN(n106) );
  NAND2_X1 U404 ( .A1(B[10]), .A2(A[10]), .ZN(n409) );
  NAND2_X1 U405 ( .A1(B[3]), .A2(A[3]), .ZN(n229) );
  NAND2_X1 U406 ( .A1(B[7]), .A2(A[7]), .ZN(n98) );
  NAND2_X1 U407 ( .A1(B[11]), .A2(A[11]), .ZN(n410) );
  NAND2_X1 U408 ( .A1(n348), .A2(n357), .ZN(n355) );
  AND2_X1 U409 ( .A1(n357), .A2(n348), .ZN(n70) );
  NAND2_X1 U410 ( .A1(B[49]), .A2(A[49]), .ZN(net495938) );
  XNOR2_X1 U411 ( .A(n188), .B(n190), .ZN(SUM[54]) );
  OAI21_X1 U412 ( .B1(n191), .B2(n511), .A(n177), .ZN(n188) );
  OAI21_X1 U413 ( .B1(n542), .B2(n1), .A(n374), .ZN(n396) );
  INV_X1 U414 ( .A(n399), .ZN(n542) );
  INV_X1 U415 ( .A(n169), .ZN(n475) );
  NAND2_X1 U416 ( .A1(B[22]), .A2(A[22]), .ZN(n325) );
  OR2_X1 U417 ( .A1(B[22]), .A2(A[22]), .ZN(n326) );
  XNOR2_X1 U418 ( .A(n33), .B(n42), .ZN(SUM[27]) );
  AOI21_X1 U419 ( .B1(n315), .B2(n12), .A(n9), .ZN(n42) );
  XNOR2_X1 U420 ( .A(n353), .B(n354), .ZN(SUM[19]) );
  OAI21_X1 U421 ( .B1(n70), .B2(n485), .A(n349), .ZN(n354) );
  AND2_X1 U422 ( .A1(B[55]), .A2(A[55]), .ZN(n86) );
  OAI211_X1 U423 ( .C1(n483), .C2(n283), .A(n341), .B(n342), .ZN(n357) );
  NAND2_X1 U424 ( .A1(n342), .A2(n348), .ZN(n359) );
  AND2_X1 U425 ( .A1(n342), .A2(n341), .ZN(n5) );
  NAND2_X1 U426 ( .A1(A[17]), .A2(B[17]), .ZN(n348) );
  NAND2_X1 U427 ( .A1(net496113), .A2(n522), .ZN(net496120) );
  INV_X1 U428 ( .A(n277), .ZN(n526) );
  OAI211_X1 U429 ( .C1(n14), .C2(n277), .A(n530), .B(n279), .ZN(n276) );
  XNOR2_X1 U430 ( .A(n22), .B(n320), .ZN(SUM[24]) );
  AOI21_X1 U431 ( .B1(n314), .B2(n319), .A(n536), .ZN(n317) );
  OAI21_X1 U432 ( .B1(n446), .B2(n277), .A(n322), .ZN(n22) );
  XNOR2_X1 U433 ( .A(net538392), .B(n255), .ZN(SUM[32]) );
  INV_X1 U434 ( .A(net538392), .ZN(n478) );
  NAND2_X1 U435 ( .A1(B[63]), .A2(A[63]), .ZN(n123) );
  NOR2_X1 U436 ( .A1(n493), .A2(n451), .ZN(net495987) );
  AND2_X1 U437 ( .A1(A[47]), .A2(B[47]), .ZN(net534711) );
  AND2_X1 U438 ( .A1(n338), .A2(n339), .ZN(n7) );
  AND2_X1 U439 ( .A1(n338), .A2(n339), .ZN(n334) );
  NAND2_X1 U440 ( .A1(net537887), .A2(n241), .ZN(n65) );
  XNOR2_X1 U441 ( .A(n211), .B(n67), .ZN(SUM[42]) );
  AOI21_X1 U442 ( .B1(n31), .B2(net495943), .A(n514), .ZN(n30) );
  INV_X1 U443 ( .A(net495943), .ZN(n515) );
  NAND2_X1 U444 ( .A1(B[53]), .A2(A[53]), .ZN(n177) );
  AOI21_X1 U445 ( .B1(n140), .B2(n141), .A(n504), .ZN(n139) );
  NOR2_X1 U446 ( .A1(n503), .A2(n505), .ZN(n140) );
  XNOR2_X1 U447 ( .A(n61), .B(n299), .ZN(SUM[29]) );
  OAI211_X1 U448 ( .C1(n516), .C2(net495937), .A(net495938), .B(net495939), 
        .ZN(net495933) );
  OAI21_X1 U449 ( .B1(n515), .B2(net538259), .A(net495937), .ZN(net538261) );
  INV_X1 U450 ( .A(net495937), .ZN(n514) );
  NAND2_X1 U451 ( .A1(n202), .A2(n203), .ZN(n201) );
  OAI21_X1 U452 ( .B1(n58), .B2(n484), .A(n362), .ZN(n360) );
  NAND2_X1 U453 ( .A1(net496035), .A2(n441), .ZN(n214) );
  NAND2_X1 U454 ( .A1(n205), .A2(n206), .ZN(n204) );
  XNOR2_X1 U455 ( .A(n215), .B(net496057), .ZN(SUM[40]) );
  NAND2_X1 U456 ( .A1(n181), .A2(n178), .ZN(n190) );
  OAI211_X1 U457 ( .C1(n482), .C2(n362), .A(n348), .B(n349), .ZN(n345) );
  INV_X1 U458 ( .A(n342), .ZN(n482) );
  OAI21_X1 U459 ( .B1(n496), .B2(n470), .A(n206), .ZN(n68) );
  INV_X1 U460 ( .A(net496057), .ZN(n470) );
  XNOR2_X1 U461 ( .A(n214), .B(n68), .ZN(SUM[41]) );
  XNOR2_X1 U462 ( .A(net538261), .B(net495961), .ZN(SUM[49]) );
  NAND2_X1 U463 ( .A1(n124), .A2(n127), .ZN(n126) );
  INV_X1 U464 ( .A(n132), .ZN(n473) );
  INV_X1 U465 ( .A(n25), .ZN(n476) );
  XNOR2_X1 U466 ( .A(n25), .B(n195), .ZN(SUM[52]) );
  XNOR2_X1 U467 ( .A(n439), .B(n303), .ZN(SUM[28]) );
  OAI21_X1 U468 ( .B1(n292), .B2(n534), .A(n265), .ZN(n62) );
  NAND2_X1 U469 ( .A1(B[60]), .A2(A[60]), .ZN(n120) );
  NAND2_X1 U470 ( .A1(n449), .A2(n243), .ZN(net495983) );
  OAI21_X1 U471 ( .B1(n232), .B2(n491), .A(n220), .ZN(n231) );
  AOI21_X1 U472 ( .B1(n521), .B2(n243), .A(n40), .ZN(n241) );
  OAI21_X1 U473 ( .B1(n497), .B2(n469), .A(n441), .ZN(n67) );
  OAI21_X1 U474 ( .B1(n469), .B2(n497), .A(n441), .ZN(n210) );
  NAND2_X1 U475 ( .A1(A[39]), .A2(B[39]), .ZN(net495986) );
  OAI21_X1 U476 ( .B1(n494), .B2(net538106), .A(net495992), .ZN(net537211) );
  XNOR2_X1 U477 ( .A(net537211), .B(n199), .ZN(SUM[46]) );
  XNOR2_X1 U478 ( .A(n133), .B(n132), .ZN(SUM[61]) );
  OAI21_X1 U479 ( .B1(n474), .B2(n506), .A(n120), .ZN(n132) );
  NAND2_X1 U480 ( .A1(n210), .A2(net496036), .ZN(n209) );
  NAND2_X1 U481 ( .A1(n153), .A2(n147), .ZN(n162) );
  INV_X1 U482 ( .A(n153), .ZN(n505) );
  XNOR2_X1 U483 ( .A(n394), .B(n393), .ZN(SUM[15]) );
  XNOR2_X1 U484 ( .A(n397), .B(n396), .ZN(SUM[14]) );
  INV_X1 U485 ( .A(n396), .ZN(n541) );
  NOR2_X1 U486 ( .A1(n514), .A2(n515), .ZN(net495965) );
  XNOR2_X1 U487 ( .A(net496010), .B(n198), .ZN(SUM[47]) );
  OAI21_X1 U488 ( .B1(n480), .B2(n533), .A(n264), .ZN(n61) );
  INV_X1 U489 ( .A(n439), .ZN(n480) );
  AOI21_X1 U490 ( .B1(n478), .B2(net496114), .A(n486), .ZN(net538497) );
  OAI221_X1 U491 ( .B1(n323), .B2(n324), .C1(n554), .C2(n525), .A(n335), .ZN(
        n280) );
  INV_X1 U492 ( .A(A[22]), .ZN(n525) );
  XNOR2_X1 U493 ( .A(n360), .B(n359), .ZN(SUM[17]) );
  NAND2_X1 U494 ( .A1(n152), .A2(n146), .ZN(n165) );
  INV_X1 U495 ( .A(n152), .ZN(n502) );
  NAND2_X1 U496 ( .A1(B[57]), .A2(A[57]), .ZN(n146) );
  OR2_X1 U497 ( .A1(B[57]), .A2(A[57]), .ZN(n152) );
  AND2_X1 U498 ( .A1(net496030), .A2(n47), .ZN(n21) );
  NAND2_X1 U499 ( .A1(net496030), .A2(n47), .ZN(net495980) );
  NAND2_X1 U500 ( .A1(n118), .A2(n128), .ZN(n127) );
  XNOR2_X1 U501 ( .A(n129), .B(n128), .ZN(SUM[62]) );
  AOI21_X1 U502 ( .B1(n302), .B2(n269), .A(n532), .ZN(n292) );
  OAI21_X1 U503 ( .B1(n481), .B2(n274), .A(n275), .ZN(n302) );
  OAI21_X1 U504 ( .B1(n24), .B2(n537), .A(n312), .ZN(n81) );
  XNOR2_X1 U505 ( .A(n24), .B(n84), .ZN(SUM[25]) );
  INV_X1 U506 ( .A(n22), .ZN(n481) );
  AOI21_X1 U507 ( .B1(n319), .B2(n314), .A(n536), .ZN(n24) );
  INV_X1 U508 ( .A(net537810), .ZN(n477) );
  NAND2_X1 U509 ( .A1(n182), .A2(n183), .ZN(n194) );
  NAND4_X1 U510 ( .A1(n183), .A2(n184), .A3(n181), .A4(n185), .ZN(n170) );
  INV_X1 U511 ( .A(n185), .ZN(n512) );
  OAI21_X1 U512 ( .B1(net538497), .B2(n247), .A(n248), .ZN(n246) );
  OR2_X1 U513 ( .A1(A[30]), .A2(B[30]), .ZN(n32) );
  NAND2_X1 U514 ( .A1(B[30]), .A2(A[30]), .ZN(n266) );
  NAND2_X1 U515 ( .A1(n237), .A2(n219), .ZN(n239) );
  INV_X1 U516 ( .A(n243), .ZN(n487) );
  NAND2_X1 U517 ( .A1(B[59]), .A2(A[59]), .ZN(n143) );
  XNOR2_X1 U518 ( .A(n191), .B(n192), .ZN(SUM[53]) );
  NOR2_X1 U519 ( .A1(n510), .A2(n511), .ZN(n192) );
  NAND2_X1 U520 ( .A1(A[14]), .A2(B[14]), .ZN(n369) );
  AND3_X1 U521 ( .A1(net496003), .A2(net495996), .A3(n10), .ZN(net538867) );
  AND4_X1 U522 ( .A1(net495996), .A2(net496003), .A3(n10), .A4(n489), .ZN(
        net495999) );
  AOI21_X1 U523 ( .B1(n53), .B2(n326), .A(n527), .ZN(n330) );
  XNOR2_X1 U524 ( .A(n442), .B(n333), .ZN(SUM[22]) );
  NAND2_X1 U525 ( .A1(n329), .A2(n328), .ZN(n338) );
  NAND2_X1 U526 ( .A1(B[19]), .A2(n438), .ZN(n282) );
  AND2_X1 U527 ( .A1(B[26]), .A2(n453), .ZN(n9) );
  OR2_X1 U528 ( .A1(B[26]), .A2(n453), .ZN(n12) );
  NAND2_X1 U529 ( .A1(A[26]), .A2(B[26]), .ZN(n52) );
  XNOR2_X1 U530 ( .A(net538259), .B(net495965), .ZN(SUM[48]) );
  NAND2_X1 U531 ( .A1(B[48]), .A2(A[48]), .ZN(net495937) );
  NAND4_X1 U532 ( .A1(n151), .A2(n152), .A3(n153), .A4(n150), .ZN(n137) );
  NAND2_X1 U533 ( .A1(n143), .A2(n150), .ZN(n158) );
  INV_X1 U534 ( .A(n150), .ZN(n503) );
  NAND2_X1 U535 ( .A1(n83), .A2(n433), .ZN(n279) );
  OAI21_X1 U536 ( .B1(n446), .B2(n277), .A(n322), .ZN(n319) );
  AOI21_X1 U537 ( .B1(n280), .B2(n83), .A(n27), .ZN(n322) );
  INV_X1 U538 ( .A(n213), .ZN(n469) );
  OAI221_X1 U539 ( .B1(n8), .B2(n23), .C1(n434), .C2(n487), .A(n522), .ZN(n216) );
  INV_X1 U540 ( .A(n38), .ZN(n521) );
  OAI22_X1 U541 ( .A1(B[35]), .A2(A[35]), .B1(B[34]), .B2(A[34]), .ZN(n38) );
  AND2_X1 U542 ( .A1(A[35]), .A2(B[35]), .ZN(n40) );
  OAI21_X1 U543 ( .B1(n471), .B2(n505), .A(n147), .ZN(n159) );
  AOI21_X1 U544 ( .B1(n173), .B2(n174), .A(n86), .ZN(n172) );
  XNOR2_X1 U546 ( .A(n62), .B(n291), .ZN(SUM[30]) );
  NAND2_X1 U547 ( .A1(n62), .A2(n32), .ZN(n290) );
  INV_X1 U548 ( .A(net495977), .ZN(n495) );
  XNOR2_X1 U549 ( .A(net496026), .B(n460), .ZN(SUM[44]) );
  NAND2_X1 U550 ( .A1(net496023), .A2(net496001), .ZN(net496022) );
  OAI21_X1 U551 ( .B1(n470), .B2(net495980), .A(net495977), .ZN(net496023) );
  NAND2_X1 U552 ( .A1(A[43]), .A2(B[43]), .ZN(n202) );
  AND2_X1 U553 ( .A1(net495985), .A2(net495986), .ZN(net495978) );
  AND4_X1 U554 ( .A1(net496008), .A2(n452), .A3(net496007), .A4(net496005), 
        .ZN(net535392) );
  AOI21_X1 U555 ( .B1(n239), .B2(n452), .A(n498), .ZN(n60) );
  AOI21_X1 U556 ( .B1(n235), .B2(n452), .A(n498), .ZN(n232) );
  NAND2_X1 U557 ( .A1(net495985), .A2(net495986), .ZN(n72) );
  AND2_X1 U558 ( .A1(net496006), .A2(net496005), .ZN(n217) );
  INV_X1 U559 ( .A(net496006), .ZN(n499) );
  OAI21_X1 U560 ( .B1(n306), .B2(n305), .A(n74), .ZN(n19) );
  OAI21_X1 U561 ( .B1(n305), .B2(n306), .A(n74), .ZN(n275) );
  NOR2_X1 U562 ( .A1(n512), .A2(n86), .ZN(n187) );
  AOI21_X1 U563 ( .B1(n259), .B2(n260), .A(n535), .ZN(n2) );
  AOI21_X1 U564 ( .B1(n259), .B2(n260), .A(n535), .ZN(n258) );
  XNOR2_X1 U565 ( .A(n457), .B(n165), .ZN(SUM[57]) );
  OAI21_X1 U566 ( .B1(n472), .B2(n502), .A(n146), .ZN(n161) );
  XNOR2_X1 U567 ( .A(n50), .B(net495948), .ZN(SUM[51]) );
  OAI21_X1 U568 ( .B1(n30), .B2(n516), .A(net495938), .ZN(net537810) );
  OAI21_X1 U569 ( .B1(n137), .B2(n475), .A(n139), .ZN(n135) );
  XNOR2_X1 U570 ( .A(n475), .B(n167), .ZN(SUM[56]) );
  OAI21_X1 U572 ( .B1(n501), .B2(n475), .A(n145), .ZN(n164) );
  OAI21_X1 U573 ( .B1(net495929), .B2(net538259), .A(n436), .ZN(n25) );
  OAI21_X1 U574 ( .B1(net495929), .B2(net538259), .A(n196), .ZN(n182) );
  NAND2_X1 U575 ( .A1(net495942), .A2(n49), .ZN(net495948) );
  NAND4_X1 U576 ( .A1(net495942), .A2(net495944), .A3(net495945), .A4(
        net495943), .ZN(net495929) );
  OAI21_X1 U577 ( .B1(n170), .B2(n476), .A(n172), .ZN(n169) );
  NOR2_X1 U578 ( .A1(n451), .A2(net534711), .ZN(net496010) );
  INV_X1 U579 ( .A(n164), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n187), .B(n186), .ZN(SUM[55]) );
  AOI21_X1 U583 ( .B1(net495932), .B2(net495933), .A(n517), .ZN(n196) );
  NAND2_X1 U584 ( .A1(B[51]), .A2(A[51]), .ZN(n49) );
  XNOR2_X1 U585 ( .A(n161), .B(n162), .ZN(SUM[58]) );
  XNOR2_X1 U586 ( .A(n159), .B(n158), .ZN(SUM[59]) );
  INV_X1 U587 ( .A(n161), .ZN(n471) );
  AOI21_X1 U588 ( .B1(n181), .B2(n188), .A(n513), .ZN(n186) );
endmodule


module RCA_NBIT64_10 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_10_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), 
        .SUM({Co, S}) );
endmodule


module RCA_NBIT64_9_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net491513, net491511, net491508, net491504, net491498, net491497,
         net491492, net491473, net491468, net491439, net538269, net538534,
         net538738, net491462, net491461, net491458, net491455, net491452,
         net491447, net491445, net491456, net491478, net491457, net491451,
         net538270, net534682, net491502, net491493, net491491, net491488,
         net491487, net491486, net491483, net491482, net491481, net491480,
         net491479, net491475, net491494, n1, n8, n9, n10, n12, n13, n14, n16,
         n17, n19, n20, n21, n22, n24, n25, n26, n30, n35, n37, n38, n40, n41,
         n42, n44, n45, n46, n49, n50, n54, n55, n56, n57, n58, n61, n64, n65,
         n66, n67, n68, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n102, n103, n104, n105, n107, n108, n109, n110, n111,
         n112, n115, n116, n119, n120, n121, n122, n124, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n137, n138, n139, n142,
         n143, n144, n145, n146, n148, n149, n150, n151, n152, n154, n156,
         n157, n159, n160, n161, n162, n163, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n175, n176, n177, n178, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n192, n193, n194,
         n195, n196, n197, n200, n202, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n222, n223, n225,
         n227, n228, n229, n230, n231, n232, n233, n236, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n253,
         n254, n255, n256, n257, n258, n260, n262, n263, n264, n267, n268,
         n270, n272, n274, n275, n276, n277, n280, n281, n282, n283, n284,
         n285, n286, n288, n289, n291, n293, n294, n295, n296, n297, n298,
         n300, n301, n302, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n318, n319, n320, n321, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n337, n338, n340, n342,
         n343, n344, n345, n346, n348, n349, n350, n351, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n369, n370, n371, n373, n374, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n398, n400, n401, n402, n403, n405,
         n406, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n423, n424, n425, n426, n427, n428, n429,
         n431, n433, n434, n435, n436, n437, n440, n441, n442, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n476, n477, n478, n479, n481, n482,
         n483, n484, n485, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614;

  OR2_X2 U10 ( .A1(B[42]), .A2(A[42]), .ZN(n194) );
  OR2_X2 U22 ( .A1(B[44]), .A2(A[44]), .ZN(n184) );
  OR2_X2 U51 ( .A1(B[50]), .A2(A[50]), .ZN(net491491) );
  NAND3_X1 U57 ( .A1(n305), .A2(n304), .A3(n306), .ZN(n295) );
  OR2_X2 U59 ( .A1(B[40]), .A2(A[40]), .ZN(n192) );
  NAND3_X1 U67 ( .A1(n394), .A2(n393), .A3(n384), .ZN(n354) );
  NAND3_X1 U68 ( .A1(n246), .A2(n240), .A3(n247), .ZN(n64) );
  NAND3_X1 U69 ( .A1(n327), .A2(n326), .A3(n406), .ZN(n318) );
  NAND3_X1 U74 ( .A1(n380), .A2(n381), .A3(n382), .ZN(n312) );
  NAND3_X1 U76 ( .A1(n280), .A2(n284), .A3(n286), .ZN(n170) );
  OR2_X2 U145 ( .A1(B[30]), .A2(A[30]), .ZN(n333) );
  NAND3_X1 U169 ( .A1(n495), .A2(n242), .A3(n19), .ZN(n236) );
  OR2_X2 U171 ( .A1(A[38]), .A2(B[38]), .ZN(n242) );
  XOR2_X1 U234 ( .A(n120), .B(n121), .Z(SUM[63]) );
  OR2_X2 U344 ( .A1(A[36]), .A2(B[36]), .ZN(n248) );
  NAND3_X1 U522 ( .A1(n195), .A2(n184), .A3(n507), .ZN(n206) );
  NAND3_X1 U524 ( .A1(n193), .A2(n213), .A3(n194), .ZN(n212) );
  NAND3_X1 U533 ( .A1(n493), .A2(n242), .A3(n243), .ZN(n240) );
  NAND3_X1 U545 ( .A1(n276), .A2(n13), .A3(n277), .ZN(n274) );
  NAND3_X1 U554 ( .A1(n309), .A2(n492), .A3(n310), .ZN(n304) );
  NAND3_X1 U555 ( .A1(n311), .A2(n312), .A3(n50), .ZN(n310) );
  NAND3_X1 U556 ( .A1(n320), .A2(n50), .A3(n321), .ZN(n294) );
  NAND3_X1 U557 ( .A1(n326), .A2(n327), .A3(n500), .ZN(n325) );
  NAND3_X1 U569 ( .A1(n377), .A2(n378), .A3(n364), .ZN(n371) );
  NAND3_X1 U570 ( .A1(n385), .A2(n384), .A3(n383), .ZN(n377) );
  NAND3_X1 U574 ( .A1(n389), .A2(n390), .A3(n313), .ZN(n382) );
  NAND3_X1 U580 ( .A1(n389), .A2(n329), .A3(n384), .ZN(n400) );
  NAND3_X1 U585 ( .A1(n405), .A2(n319), .A3(n318), .ZN(n384) );
  NAND3_X1 U586 ( .A1(n326), .A2(n497), .A3(n411), .ZN(n405) );
  NAND3_X1 U598 ( .A1(n464), .A2(n465), .A3(n466), .ZN(n463) );
  NAND3_X1 U599 ( .A1(n467), .A2(n85), .A3(n468), .ZN(n464) );
  OR2_X2 U40 ( .A1(A[25]), .A2(B[25]), .ZN(n361) );
  OR2_X2 U128 ( .A1(B[52]), .A2(A[52]), .ZN(net491456) );
  OR2_X2 U138 ( .A1(B[54]), .A2(A[54]), .ZN(net491455) );
  OR2_X2 U361 ( .A1(B[41]), .A2(A[41]), .ZN(n193) );
  OR2_X2 U365 ( .A1(B[57]), .A2(A[57]), .ZN(n144) );
  OR2_X2 U392 ( .A1(B[58]), .A2(A[58]), .ZN(n142) );
  CLKBUF_X1 U2 ( .A(A[47]), .Z(n489) );
  AND2_X1 U3 ( .A1(n423), .A2(n408), .ZN(n420) );
  INV_X1 U4 ( .A(n300), .ZN(n582) );
  OR2_X1 U5 ( .A1(n580), .A2(n581), .ZN(n508) );
  OR2_X1 U6 ( .A1(A[33]), .A2(B[33]), .ZN(n288) );
  NOR2_X1 U7 ( .A1(B[32]), .A2(A[32]), .ZN(n74) );
  OR2_X1 U8 ( .A1(B[49]), .A2(A[49]), .ZN(net491493) );
  AND2_X1 U9 ( .A1(n481), .A2(n413), .ZN(SUM[0]) );
  AND2_X1 U11 ( .A1(n501), .A2(n361), .ZN(n490) );
  AND2_X1 U12 ( .A1(n369), .A2(n359), .ZN(n491) );
  CLKBUF_X1 U13 ( .A(n308), .Z(n492) );
  OR2_X2 U14 ( .A1(A[37]), .A2(B[37]), .ZN(n493) );
  OR2_X1 U15 ( .A1(B[37]), .A2(A[37]), .ZN(n241) );
  OR2_X1 U16 ( .A1(B[23]), .A2(A[23]), .ZN(n311) );
  CLKBUF_X1 U17 ( .A(n166), .Z(n494) );
  OR2_X1 U18 ( .A1(A[39]), .A2(B[39]), .ZN(n495) );
  OR2_X1 U19 ( .A1(A[39]), .A2(B[39]), .ZN(n238) );
  OR2_X2 U20 ( .A1(B[18]), .A2(A[18]), .ZN(n326) );
  AOI21_X1 U21 ( .B1(n297), .B2(n298), .A(n76), .ZN(n496) );
  CLKBUF_X1 U23 ( .A(n337), .Z(n497) );
  NAND2_X1 U24 ( .A1(n67), .A2(n68), .ZN(n498) );
  NAND2_X1 U25 ( .A1(n371), .A2(n490), .ZN(n370) );
  CLKBUF_X1 U26 ( .A(n437), .Z(n499) );
  OR2_X1 U27 ( .A1(A[15]), .A2(B[15]), .ZN(n437) );
  OR2_X1 U28 ( .A1(B[56]), .A2(A[56]), .ZN(n143) );
  CLKBUF_X1 U29 ( .A(n328), .Z(n500) );
  OR2_X2 U30 ( .A1(A[22]), .A2(B[22]), .ZN(n313) );
  OR2_X1 U31 ( .A1(B[26]), .A2(A[26]), .ZN(n501) );
  OR2_X1 U32 ( .A1(B[26]), .A2(A[26]), .ZN(n362) );
  NAND3_X1 U33 ( .A1(n305), .A2(n304), .A3(n306), .ZN(n502) );
  AND2_X1 U34 ( .A1(n409), .A2(n330), .ZN(n421) );
  OR2_X2 U35 ( .A1(A[17]), .A2(B[17]), .ZN(n330) );
  OR2_X1 U36 ( .A1(A[47]), .A2(B[47]), .ZN(n503) );
  CLKBUF_X1 U37 ( .A(n301), .Z(n504) );
  NAND3_X1 U38 ( .A1(n493), .A2(n242), .A3(n243), .ZN(n505) );
  NAND2_X1 U39 ( .A1(n370), .A2(n491), .ZN(n366) );
  INV_X1 U41 ( .A(n13), .ZN(n506) );
  NAND2_X1 U42 ( .A1(n211), .A2(n212), .ZN(n507) );
  OR2_X1 U43 ( .A1(B[43]), .A2(A[43]), .ZN(n195) );
  XNOR2_X1 U44 ( .A(n340), .B(n508), .ZN(SUM[30]) );
  OR2_X2 U45 ( .A1(B[53]), .A2(A[53]), .ZN(net491457) );
  OAI211_X1 U46 ( .C1(n574), .C2(n281), .A(n282), .B(n283), .ZN(n509) );
  OAI21_X1 U47 ( .B1(n568), .B2(n30), .A(net491451), .ZN(n510) );
  NOR2_X1 U48 ( .A1(A[34]), .A2(B[34]), .ZN(n190) );
  OR2_X1 U49 ( .A1(B[35]), .A2(A[35]), .ZN(n189) );
  NOR2_X1 U50 ( .A1(B[55]), .A2(A[55]), .ZN(n511) );
  NAND3_X1 U52 ( .A1(n509), .A2(n284), .A3(n286), .ZN(n512) );
  XNOR2_X1 U53 ( .A(n338), .B(n513), .ZN(SUM[31]) );
  NOR2_X1 U54 ( .A1(n76), .A2(n45), .ZN(n513) );
  CLKBUF_X1 U55 ( .A(n227), .Z(n514) );
  AND2_X1 U56 ( .A1(A[46]), .A2(B[46]), .ZN(n515) );
  OR2_X1 U58 ( .A1(B[46]), .A2(A[46]), .ZN(n177) );
  NOR2_X1 U60 ( .A1(B[59]), .A2(A[59]), .ZN(n516) );
  XOR2_X1 U61 ( .A(n532), .B(n517), .Z(SUM[45]) );
  OR2_X1 U62 ( .A1(n544), .A2(n546), .ZN(n517) );
  XNOR2_X1 U63 ( .A(n9), .B(n518), .ZN(SUM[28]) );
  OR2_X1 U64 ( .A1(n582), .A2(n583), .ZN(n518) );
  XNOR2_X1 U65 ( .A(n17), .B(n519), .ZN(SUM[34]) );
  OR2_X1 U66 ( .A1(n77), .A2(n190), .ZN(n519) );
  OAI211_X1 U70 ( .C1(n293), .C2(n294), .A(n295), .B(n296), .ZN(n187) );
  NOR2_X1 U71 ( .A1(n585), .A2(n584), .ZN(n376) );
  NOR2_X1 U72 ( .A1(n552), .A2(n553), .ZN(n275) );
  XOR2_X1 U73 ( .A(n520), .B(n398), .Z(SUM[22]) );
  NOR2_X1 U75 ( .A1(n593), .A2(n592), .ZN(n520) );
  AOI21_X1 U77 ( .B1(n187), .B2(n575), .A(n576), .ZN(n26) );
  OAI21_X1 U78 ( .B1(n163), .B2(n541), .A(n72), .ZN(n162) );
  AOI21_X1 U79 ( .B1(n494), .B2(n167), .A(n168), .ZN(n163) );
  NAND2_X1 U80 ( .A1(n536), .A2(n169), .ZN(n167) );
  NAND2_X1 U81 ( .A1(n14), .A2(n166), .ZN(n218) );
  INV_X1 U82 ( .A(net491475), .ZN(n530) );
  INV_X1 U83 ( .A(A[26]), .ZN(n586) );
  AND2_X1 U84 ( .A1(n189), .A2(n575), .ZN(n277) );
  INV_X1 U85 ( .A(n236), .ZN(n536) );
  AND3_X1 U86 ( .A1(n276), .A2(n13), .A3(n277), .ZN(n1) );
  OAI21_X1 U87 ( .B1(n610), .B2(n449), .A(n446), .ZN(n88) );
  NOR2_X1 U88 ( .A1(n442), .A2(n599), .ZN(n425) );
  INV_X1 U89 ( .A(n444), .ZN(n599) );
  AOI21_X1 U90 ( .B1(n445), .B2(n446), .A(n447), .ZN(n442) );
  NAND2_X1 U91 ( .A1(n602), .A2(n448), .ZN(n445) );
  NAND2_X1 U92 ( .A1(n461), .A2(n444), .ZN(n459) );
  NAND2_X1 U93 ( .A1(n598), .A2(n88), .ZN(n461) );
  INV_X1 U94 ( .A(n447), .ZN(n598) );
  INV_X1 U95 ( .A(n448), .ZN(n610) );
  INV_X1 U96 ( .A(n449), .ZN(n602) );
  NOR2_X1 U97 ( .A1(n105), .A2(n558), .ZN(SUM[64]) );
  AND2_X1 U98 ( .A1(n171), .A2(n284), .ZN(n66) );
  NAND2_X1 U99 ( .A1(n214), .A2(n193), .ZN(n228) );
  AOI21_X1 U100 ( .B1(n119), .B2(n122), .A(n559), .ZN(n120) );
  NAND2_X1 U101 ( .A1(n111), .A2(n107), .ZN(n121) );
  INV_X1 U102 ( .A(n112), .ZN(n559) );
  OAI211_X1 U103 ( .C1(n577), .C2(n300), .A(n504), .B(n302), .ZN(n298) );
  INV_X1 U104 ( .A(n307), .ZN(n577) );
  NAND2_X1 U105 ( .A1(n115), .A2(n126), .ZN(n128) );
  NAND2_X1 U106 ( .A1(n194), .A2(n217), .ZN(n225) );
  NAND2_X1 U107 ( .A1(net491455), .A2(net491452), .ZN(net491468) );
  NAND2_X1 U108 ( .A1(n142), .A2(n139), .ZN(n154) );
  XNOR2_X1 U109 ( .A(n374), .B(n373), .ZN(SUM[26]) );
  XNOR2_X1 U110 ( .A(n387), .B(n386), .ZN(SUM[24]) );
  NAND2_X1 U111 ( .A1(n365), .A2(n364), .ZN(n386) );
  NAND2_X1 U112 ( .A1(n311), .A2(n312), .ZN(n388) );
  OAI211_X1 U113 ( .C1(n589), .C2(n392), .A(n391), .B(n400), .ZN(n398) );
  XNOR2_X1 U114 ( .A(n267), .B(n268), .ZN(SUM[37]) );
  NOR2_X1 U115 ( .A1(n537), .A2(n538), .ZN(n268) );
  INV_X1 U116 ( .A(n493), .ZN(n538) );
  OAI211_X1 U117 ( .C1(n557), .C2(n137), .A(n138), .B(n139), .ZN(n135) );
  XOR2_X1 U118 ( .A(n218), .B(n521), .Z(SUM[40]) );
  AND2_X1 U119 ( .A1(n192), .A2(n215), .ZN(n521) );
  XNOR2_X1 U120 ( .A(n395), .B(n396), .ZN(SUM[23]) );
  NOR2_X1 U121 ( .A1(n591), .A2(n71), .ZN(n396) );
  AOI21_X1 U122 ( .B1(n313), .B2(n398), .A(n592), .ZN(n395) );
  INV_X1 U123 ( .A(n380), .ZN(n591) );
  XNOR2_X1 U124 ( .A(n415), .B(n414), .ZN(SUM[19]) );
  NAND2_X1 U125 ( .A1(n319), .A2(n327), .ZN(n414) );
  NAND2_X1 U126 ( .A1(n417), .A2(n416), .ZN(n415) );
  OAI211_X1 U127 ( .C1(n568), .C2(n38), .A(net491451), .B(net491452), .ZN(
        net491447) );
  AOI21_X1 U129 ( .B1(net491456), .B2(net491475), .A(n563), .ZN(n30) );
  INV_X1 U130 ( .A(n38), .ZN(n563) );
  NAND2_X1 U131 ( .A1(n493), .A2(n248), .ZN(n263) );
  AOI21_X1 U132 ( .B1(n552), .B2(n493), .A(n537), .ZN(n264) );
  NAND2_X1 U133 ( .A1(n181), .A2(n184), .ZN(n209) );
  NAND2_X1 U134 ( .A1(n38), .A2(net491456), .ZN(net491478) );
  NAND2_X1 U135 ( .A1(n138), .A2(n144), .ZN(n157) );
  NOR2_X1 U136 ( .A1(n168), .A2(n186), .ZN(n172) );
  NAND4_X1 U137 ( .A1(n536), .A2(n188), .A3(n189), .A4(n13), .ZN(n186) );
  OAI211_X1 U139 ( .C1(n207), .C2(n549), .A(n206), .B(n181), .ZN(n35) );
  INV_X1 U140 ( .A(n184), .ZN(n549) );
  NOR3_X1 U141 ( .A1(n190), .A2(n574), .A3(n74), .ZN(n188) );
  XNOR2_X1 U142 ( .A(n366), .B(n367), .ZN(SUM[27]) );
  NAND2_X1 U143 ( .A1(n61), .A2(n360), .ZN(n367) );
  INV_X1 U144 ( .A(n139), .ZN(n555) );
  NAND2_X1 U146 ( .A1(n116), .A2(n129), .ZN(n131) );
  XNOR2_X1 U147 ( .A(n46), .B(n289), .ZN(SUM[33]) );
  NAND2_X1 U148 ( .A1(n282), .A2(n288), .ZN(n289) );
  OAI21_X1 U149 ( .B1(n524), .B2(n74), .A(n281), .ZN(n46) );
  XNOR2_X1 U150 ( .A(n122), .B(n124), .ZN(SUM[62]) );
  NAND2_X1 U151 ( .A1(n119), .A2(n112), .ZN(n124) );
  XOR2_X1 U152 ( .A(n522), .B(net491513), .Z(SUM[48]) );
  AND2_X1 U153 ( .A1(net491486), .A2(net491492), .ZN(n522) );
  XNOR2_X1 U154 ( .A(n401), .B(n402), .ZN(SUM[21]) );
  NAND2_X1 U155 ( .A1(n389), .A2(n391), .ZN(n401) );
  OAI21_X1 U156 ( .B1(n22), .B2(n587), .A(n392), .ZN(n402) );
  XNOR2_X1 U157 ( .A(n350), .B(n349), .ZN(SUM[29]) );
  NAND2_X1 U158 ( .A1(n307), .A2(n504), .ZN(n349) );
  NAND2_X1 U159 ( .A1(n342), .A2(n300), .ZN(n350) );
  XNOR2_X1 U160 ( .A(n506), .B(n291), .ZN(SUM[32]) );
  NOR2_X1 U161 ( .A1(n576), .A2(n74), .ZN(n291) );
  XNOR2_X1 U162 ( .A(n424), .B(n25), .ZN(SUM[16]) );
  NAND2_X1 U163 ( .A1(n328), .A2(n408), .ZN(n424) );
  XNOR2_X1 U164 ( .A(n257), .B(n258), .ZN(SUM[39]) );
  NOR2_X1 U165 ( .A1(n539), .A2(n540), .ZN(n258) );
  XNOR2_X1 U166 ( .A(n22), .B(n403), .ZN(SUM[20]) );
  NOR2_X1 U167 ( .A1(n588), .A2(n587), .ZN(n403) );
  INV_X1 U168 ( .A(n392), .ZN(n588) );
  XNOR2_X1 U170 ( .A(n57), .B(n419), .ZN(SUM[18]) );
  NAND2_X1 U172 ( .A1(n326), .A2(n416), .ZN(n419) );
  OAI21_X1 U173 ( .B1(n420), .B2(n534), .A(n409), .ZN(n57) );
  XNOR2_X1 U174 ( .A(n222), .B(n58), .ZN(SUM[43]) );
  AOI21_X1 U175 ( .B1(n223), .B2(n194), .A(n542), .ZN(n222) );
  INV_X1 U176 ( .A(n217), .ZN(n542) );
  NAND4_X1 U177 ( .A1(n195), .A2(n193), .A3(n194), .A4(n192), .ZN(n168) );
  NAND2_X1 U178 ( .A1(net538270), .A2(net491481), .ZN(net491475) );
  AOI21_X1 U179 ( .B1(net491482), .B2(net491483), .A(net534682), .ZN(net491481) );
  INV_X1 U180 ( .A(net491513), .ZN(n531) );
  NAND2_X1 U181 ( .A1(net491491), .A2(net491488), .ZN(net491504) );
  OAI21_X1 U182 ( .B1(n527), .B2(n562), .A(n116), .ZN(n127) );
  INV_X1 U183 ( .A(net491452), .ZN(n567) );
  NAND2_X1 U184 ( .A1(n391), .A2(n392), .ZN(n390) );
  NOR2_X1 U185 ( .A1(n324), .A2(n325), .ZN(n320) );
  OAI211_X1 U186 ( .C1(n596), .C2(n433), .A(n434), .B(n435), .ZN(n429) );
  NAND4_X1 U187 ( .A1(n331), .A2(n332), .A3(n307), .A4(n333), .ZN(n293) );
  NOR3_X1 U188 ( .A1(n71), .A2(n589), .A3(n593), .ZN(n332) );
  NOR2_X1 U189 ( .A1(n594), .A2(n583), .ZN(n331) );
  INV_X1 U190 ( .A(n25), .ZN(n594) );
  AND2_X1 U191 ( .A1(n44), .A2(n12), .ZN(n306) );
  XNOR2_X1 U192 ( .A(n80), .B(n202), .ZN(SUM[46]) );
  OAI21_X1 U193 ( .B1(n532), .B2(n546), .A(n182), .ZN(n80) );
  NAND4_X1 U194 ( .A1(n219), .A2(n218), .A3(n195), .A4(n194), .ZN(n207) );
  NOR2_X1 U195 ( .A1(n543), .A2(n551), .ZN(n219) );
  INV_X1 U196 ( .A(n192), .ZN(n551) );
  XNOR2_X1 U197 ( .A(net538269), .B(net491473), .ZN(SUM[53]) );
  OAI21_X1 U198 ( .B1(n564), .B2(n530), .A(n38), .ZN(net538269) );
  INV_X1 U199 ( .A(net491456), .ZN(n564) );
  AOI21_X1 U200 ( .B1(n573), .B2(n248), .A(n552), .ZN(n272) );
  INV_X1 U201 ( .A(n171), .ZN(n573) );
  INV_X1 U202 ( .A(n288), .ZN(n574) );
  INV_X1 U203 ( .A(n329), .ZN(n587) );
  INV_X1 U204 ( .A(n389), .ZN(n589) );
  INV_X1 U205 ( .A(n182), .ZN(n544) );
  INV_X1 U206 ( .A(n330), .ZN(n534) );
  NOR2_X1 U207 ( .A1(n547), .A2(n548), .ZN(n197) );
  AOI21_X1 U208 ( .B1(n200), .B2(n177), .A(n515), .ZN(n196) );
  AND3_X1 U209 ( .A1(n405), .A2(n319), .A3(n318), .ZN(n22) );
  OAI21_X1 U210 ( .B1(n543), .B2(n533), .A(n214), .ZN(n223) );
  OAI21_X1 U211 ( .B1(n532), .B2(n546), .A(n182), .ZN(n200) );
  AND2_X1 U212 ( .A1(n185), .A2(n184), .ZN(n10) );
  AOI21_X1 U213 ( .B1(n428), .B2(n429), .A(n595), .ZN(n427) );
  AND2_X1 U214 ( .A1(n437), .A2(n436), .ZN(n428) );
  INV_X1 U215 ( .A(n313), .ZN(n593) );
  INV_X1 U216 ( .A(n185), .ZN(n546) );
  OAI21_X1 U217 ( .B1(n425), .B2(n426), .A(n24), .ZN(n25) );
  AOI21_X1 U218 ( .B1(n21), .B2(n429), .A(n595), .ZN(n24) );
  AND2_X1 U219 ( .A1(n437), .A2(n436), .ZN(n21) );
  NAND2_X1 U220 ( .A1(n244), .A2(n245), .ZN(n243) );
  INV_X1 U221 ( .A(net491455), .ZN(n566) );
  INV_X1 U222 ( .A(n142), .ZN(n556) );
  NOR2_X1 U223 ( .A1(n574), .A2(n190), .ZN(n276) );
  NOR2_X1 U224 ( .A1(n593), .A2(n71), .ZN(n385) );
  AND3_X1 U225 ( .A1(n365), .A2(n389), .A3(n329), .ZN(n383) );
  AND3_X1 U226 ( .A1(n327), .A2(n330), .A3(n500), .ZN(n411) );
  OR2_X1 U227 ( .A1(n578), .A2(n82), .ZN(n68) );
  INV_X1 U228 ( .A(n81), .ZN(n578) );
  INV_X1 U229 ( .A(n245), .ZN(n552) );
  NAND4_X1 U230 ( .A1(n313), .A2(n314), .A3(n315), .A4(n50), .ZN(n309) );
  NAND2_X1 U231 ( .A1(n318), .A2(n319), .ZN(n314) );
  NOR3_X1 U232 ( .A1(n71), .A2(n589), .A3(n587), .ZN(n315) );
  NAND2_X1 U233 ( .A1(n337), .A2(n328), .ZN(n423) );
  OAI21_X1 U235 ( .B1(n420), .B2(n534), .A(n409), .ZN(n418) );
  NAND2_X1 U236 ( .A1(n214), .A2(n215), .ZN(n213) );
  NOR2_X1 U237 ( .A1(n570), .A2(net534682), .ZN(net491498) );
  INV_X1 U238 ( .A(net491488), .ZN(n571) );
  NAND2_X1 U239 ( .A1(n238), .A2(n233), .ZN(n166) );
  INV_X1 U240 ( .A(n193), .ZN(n543) );
  INV_X1 U241 ( .A(n74), .ZN(n575) );
  INV_X1 U242 ( .A(n361), .ZN(n584) );
  INV_X1 U243 ( .A(n281), .ZN(n576) );
  INV_X1 U244 ( .A(n431), .ZN(n595) );
  AND3_X1 U245 ( .A1(n377), .A2(n364), .A3(n378), .ZN(n54) );
  INV_X1 U246 ( .A(n129), .ZN(n562) );
  INV_X1 U247 ( .A(n244), .ZN(n537) );
  INV_X1 U248 ( .A(n363), .ZN(n585) );
  NAND2_X1 U249 ( .A1(n607), .A2(n572), .ZN(n284) );
  INV_X1 U250 ( .A(n248), .ZN(n553) );
  INV_X1 U251 ( .A(net491493), .ZN(n565) );
  NAND2_X1 U252 ( .A1(n55), .A2(n379), .ZN(n378) );
  AND2_X1 U253 ( .A1(n365), .A2(n311), .ZN(n379) );
  NAND2_X1 U254 ( .A1(n8), .A2(n382), .ZN(n55) );
  AND2_X1 U255 ( .A1(n380), .A2(n381), .ZN(n8) );
  INV_X1 U256 ( .A(n305), .ZN(n583) );
  NAND2_X1 U257 ( .A1(n329), .A2(n330), .ZN(n324) );
  INV_X1 U258 ( .A(n381), .ZN(n592) );
  INV_X1 U259 ( .A(n126), .ZN(n561) );
  INV_X1 U260 ( .A(n144), .ZN(n557) );
  OR2_X1 U261 ( .A1(n353), .A2(n56), .ZN(n355) );
  NAND2_X1 U262 ( .A1(n312), .A2(n311), .ZN(n56) );
  INV_X1 U263 ( .A(n333), .ZN(n581) );
  INV_X1 U264 ( .A(n302), .ZN(n580) );
  INV_X1 U265 ( .A(net491508), .ZN(n525) );
  AND2_X1 U266 ( .A1(n241), .A2(n248), .ZN(n19) );
  INV_X1 U267 ( .A(n176), .ZN(n548) );
  INV_X1 U268 ( .A(n495), .ZN(n540) );
  INV_X1 U269 ( .A(n215), .ZN(n550) );
  AND2_X1 U270 ( .A1(n300), .A2(n301), .ZN(n82) );
  AND2_X1 U271 ( .A1(n363), .A2(n364), .ZN(n73) );
  AND2_X1 U272 ( .A1(n333), .A2(n307), .ZN(n12) );
  AND2_X1 U273 ( .A1(n305), .A2(n81), .ZN(n79) );
  INV_X1 U274 ( .A(n247), .ZN(n535) );
  XNOR2_X1 U275 ( .A(n450), .B(n451), .ZN(SUM[15]) );
  NAND2_X1 U276 ( .A1(n452), .A2(n435), .ZN(n451) );
  NAND2_X1 U277 ( .A1(n431), .A2(n499), .ZN(n450) );
  NAND2_X1 U278 ( .A1(n436), .A2(n453), .ZN(n452) );
  XNOR2_X1 U279 ( .A(n454), .B(n453), .ZN(SUM[14]) );
  NAND2_X1 U280 ( .A1(n436), .A2(n435), .ZN(n454) );
  XNOR2_X1 U281 ( .A(n457), .B(n456), .ZN(SUM[13]) );
  NAND2_X1 U282 ( .A1(n441), .A2(n434), .ZN(n457) );
  XNOR2_X1 U283 ( .A(n91), .B(n92), .ZN(SUM[7]) );
  NAND2_X1 U284 ( .A1(n95), .A2(n96), .ZN(n91) );
  NAND2_X1 U285 ( .A1(n93), .A2(n94), .ZN(n92) );
  NAND2_X1 U286 ( .A1(n97), .A2(n98), .ZN(n96) );
  XNOR2_X1 U287 ( .A(n469), .B(n470), .ZN(SUM[11]) );
  NAND2_X1 U288 ( .A1(n465), .A2(n471), .ZN(n470) );
  NAND2_X1 U289 ( .A1(n466), .A2(n462), .ZN(n469) );
  NAND2_X1 U290 ( .A1(n468), .A2(n472), .ZN(n471) );
  XNOR2_X1 U291 ( .A(n249), .B(n250), .ZN(SUM[3]) );
  OAI21_X1 U292 ( .B1(n613), .B2(n611), .A(n253), .ZN(n250) );
  NAND2_X1 U293 ( .A1(n255), .A2(n256), .ZN(n249) );
  INV_X1 U294 ( .A(n254), .ZN(n613) );
  XNOR2_X1 U295 ( .A(n412), .B(n614), .ZN(SUM[1]) );
  NAND2_X1 U296 ( .A1(n346), .A2(n345), .ZN(n412) );
  XNOR2_X1 U297 ( .A(n460), .B(n459), .ZN(SUM[12]) );
  NAND2_X1 U298 ( .A1(n440), .A2(n433), .ZN(n460) );
  XNOR2_X1 U299 ( .A(n87), .B(n88), .ZN(SUM[8]) );
  NAND2_X1 U300 ( .A1(n89), .A2(n90), .ZN(n87) );
  XNOR2_X1 U301 ( .A(n83), .B(n84), .ZN(SUM[9]) );
  NAND2_X1 U302 ( .A1(n85), .A2(n86), .ZN(n83) );
  XNOR2_X1 U303 ( .A(n146), .B(n104), .ZN(SUM[5]) );
  NAND2_X1 U304 ( .A1(n103), .A2(n102), .ZN(n146) );
  XNOR2_X1 U305 ( .A(n99), .B(n97), .ZN(SUM[6]) );
  NAND2_X1 U306 ( .A1(n98), .A2(n95), .ZN(n99) );
  XNOR2_X1 U307 ( .A(n473), .B(n472), .ZN(SUM[10]) );
  NAND2_X1 U308 ( .A1(n468), .A2(n465), .ZN(n473) );
  XNOR2_X1 U309 ( .A(n343), .B(n254), .ZN(SUM[2]) );
  NAND2_X1 U310 ( .A1(n348), .A2(n253), .ZN(n343) );
  XNOR2_X1 U311 ( .A(n160), .B(n448), .ZN(SUM[4]) );
  NAND2_X1 U312 ( .A1(n149), .A2(n148), .ZN(n160) );
  OAI21_X1 U313 ( .B1(n482), .B2(n483), .A(n256), .ZN(n448) );
  NAND2_X1 U314 ( .A1(n348), .A2(n255), .ZN(n483) );
  NOR2_X1 U315 ( .A1(n484), .A2(n485), .ZN(n482) );
  NAND2_X1 U316 ( .A1(n253), .A2(n345), .ZN(n485) );
  OAI21_X1 U317 ( .B1(n601), .B2(n600), .A(n86), .ZN(n472) );
  INV_X1 U318 ( .A(n84), .ZN(n601) );
  INV_X1 U319 ( .A(n85), .ZN(n600) );
  OAI21_X1 U320 ( .B1(n597), .B2(n596), .A(n434), .ZN(n453) );
  INV_X1 U321 ( .A(n456), .ZN(n597) );
  OAI21_X1 U322 ( .B1(n605), .B2(n610), .A(n148), .ZN(n104) );
  INV_X1 U323 ( .A(n149), .ZN(n605) );
  OAI21_X1 U324 ( .B1(n604), .B2(n603), .A(n102), .ZN(n97) );
  INV_X1 U325 ( .A(n104), .ZN(n604) );
  INV_X1 U326 ( .A(n103), .ZN(n603) );
  OAI21_X1 U327 ( .B1(n477), .B2(n478), .A(n93), .ZN(n446) );
  NAND2_X1 U328 ( .A1(n94), .A2(n95), .ZN(n478) );
  NOR2_X1 U329 ( .A1(n20), .A2(n479), .ZN(n477) );
  AND2_X1 U330 ( .A1(n102), .A2(n148), .ZN(n20) );
  NAND4_X1 U331 ( .A1(n149), .A2(n103), .A3(n98), .A4(n93), .ZN(n449) );
  NAND4_X1 U332 ( .A1(n85), .A2(n89), .A3(n468), .A4(n462), .ZN(n447) );
  AOI21_X1 U333 ( .B1(n108), .B2(n109), .A(n110), .ZN(n105) );
  NAND2_X1 U334 ( .A1(n111), .A2(n112), .ZN(n110) );
  NOR2_X1 U335 ( .A1(n560), .A2(n561), .ZN(n108) );
  OAI211_X1 U336 ( .C1(n527), .C2(n562), .A(n115), .B(n116), .ZN(n109) );
  NAND4_X1 U337 ( .A1(n440), .A2(n441), .A3(n436), .A4(n499), .ZN(n426) );
  NOR2_X1 U338 ( .A1(n612), .A2(n413), .ZN(n484) );
  INV_X1 U339 ( .A(n346), .ZN(n612) );
  NAND2_X1 U340 ( .A1(n476), .A2(n90), .ZN(n84) );
  NAND2_X1 U341 ( .A1(n88), .A2(n89), .ZN(n476) );
  NAND2_X1 U342 ( .A1(n344), .A2(n345), .ZN(n254) );
  NAND2_X1 U343 ( .A1(n346), .A2(n614), .ZN(n344) );
  NAND2_X1 U345 ( .A1(n458), .A2(n433), .ZN(n456) );
  NAND2_X1 U346 ( .A1(n459), .A2(n440), .ZN(n458) );
  NAND2_X1 U347 ( .A1(n462), .A2(n463), .ZN(n444) );
  NAND2_X1 U348 ( .A1(n86), .A2(n90), .ZN(n467) );
  INV_X1 U349 ( .A(n413), .ZN(n614) );
  INV_X1 U350 ( .A(n441), .ZN(n596) );
  NAND2_X1 U351 ( .A1(n103), .A2(n98), .ZN(n479) );
  INV_X1 U352 ( .A(n348), .ZN(n611) );
  INV_X1 U353 ( .A(n119), .ZN(n560) );
  INV_X1 U354 ( .A(n107), .ZN(n558) );
  NOR2_X1 U355 ( .A1(B[23]), .A2(A[23]), .ZN(n71) );
  NAND2_X1 U356 ( .A1(B[26]), .A2(A[26]), .ZN(n359) );
  OAI211_X1 U357 ( .C1(n534), .C2(n408), .A(n409), .B(n410), .ZN(n406) );
  OAI211_X1 U358 ( .C1(n574), .C2(n281), .A(n282), .B(n283), .ZN(n280) );
  NAND2_X1 U359 ( .A1(B[34]), .A2(A[34]), .ZN(n283) );
  NAND2_X1 U360 ( .A1(B[20]), .A2(A[20]), .ZN(n392) );
  NAND2_X1 U362 ( .A1(B[52]), .A2(A[52]), .ZN(n38) );
  NOR2_X1 U363 ( .A1(n589), .A2(n587), .ZN(n393) );
  AOI21_X1 U364 ( .B1(n606), .B2(n590), .A(n593), .ZN(n394) );
  INV_X1 U366 ( .A(B[23]), .ZN(n606) );
  NAND2_X1 U367 ( .A1(B[28]), .A2(A[28]), .ZN(n300) );
  OR2_X1 U368 ( .A1(A[14]), .A2(B[14]), .ZN(n436) );
  NAND2_X1 U369 ( .A1(B[45]), .A2(A[45]), .ZN(n182) );
  NAND2_X1 U370 ( .A1(B[41]), .A2(A[41]), .ZN(n214) );
  NAND2_X1 U371 ( .A1(A[19]), .A2(B[19]), .ZN(n319) );
  NAND2_X1 U372 ( .A1(A[14]), .A2(B[14]), .ZN(n435) );
  OR2_X1 U373 ( .A1(B[24]), .A2(A[24]), .ZN(n365) );
  OR2_X1 U374 ( .A1(B[21]), .A2(A[21]), .ZN(n389) );
  NAND2_X1 U375 ( .A1(B[33]), .A2(A[33]), .ZN(n282) );
  NAND2_X1 U376 ( .A1(B[62]), .A2(A[62]), .ZN(n112) );
  NAND2_X1 U377 ( .A1(B[40]), .A2(A[40]), .ZN(n215) );
  NAND2_X1 U378 ( .A1(B[32]), .A2(A[32]), .ZN(n281) );
  NAND2_X1 U379 ( .A1(B[58]), .A2(A[58]), .ZN(n139) );
  NAND2_X1 U380 ( .A1(B[54]), .A2(A[54]), .ZN(net491452) );
  OR2_X1 U381 ( .A1(A[29]), .A2(B[29]), .ZN(n307) );
  NAND2_X1 U382 ( .A1(B[21]), .A2(A[21]), .ZN(n391) );
  NAND2_X1 U383 ( .A1(B[24]), .A2(A[24]), .ZN(n364) );
  NAND2_X1 U384 ( .A1(B[61]), .A2(A[61]), .ZN(n115) );
  NAND2_X1 U385 ( .A1(B[50]), .A2(A[50]), .ZN(net491488) );
  OR2_X1 U386 ( .A1(A[16]), .A2(B[16]), .ZN(n328) );
  NAND2_X1 U387 ( .A1(A[16]), .A2(B[16]), .ZN(n408) );
  NAND2_X1 U388 ( .A1(B[44]), .A2(A[44]), .ZN(n181) );
  NAND2_X1 U389 ( .A1(B[57]), .A2(A[57]), .ZN(n138) );
  OR2_X1 U390 ( .A1(A[20]), .A2(B[20]), .ZN(n329) );
  NAND2_X1 U391 ( .A1(A[38]), .A2(B[38]), .ZN(n247) );
  NAND2_X1 U393 ( .A1(B[42]), .A2(A[42]), .ZN(n217) );
  OR2_X1 U394 ( .A1(B[62]), .A2(A[62]), .ZN(n119) );
  NAND2_X1 U395 ( .A1(B[49]), .A2(A[49]), .ZN(net491487) );
  OR2_X1 U396 ( .A1(A[19]), .A2(B[19]), .ZN(n327) );
  OR2_X1 U397 ( .A1(B[28]), .A2(A[28]), .ZN(n305) );
  NAND2_X1 U398 ( .A1(A[46]), .A2(B[46]), .ZN(n183) );
  NAND2_X1 U399 ( .A1(B[53]), .A2(A[53]), .ZN(net491451) );
  NAND2_X1 U400 ( .A1(A[22]), .A2(B[22]), .ZN(n381) );
  NAND2_X1 U401 ( .A1(n489), .A2(B[47]), .ZN(n176) );
  NAND2_X1 U402 ( .A1(A[39]), .A2(B[39]), .ZN(n246) );
  NAND2_X1 U403 ( .A1(B[30]), .A2(A[30]), .ZN(n302) );
  NAND2_X1 U404 ( .A1(A[36]), .A2(B[36]), .ZN(n245) );
  NAND2_X1 U405 ( .A1(B[37]), .A2(A[37]), .ZN(n244) );
  NAND2_X1 U406 ( .A1(B[63]), .A2(A[63]), .ZN(n111) );
  OR2_X1 U407 ( .A1(B[61]), .A2(A[61]), .ZN(n126) );
  OR2_X1 U408 ( .A1(B[63]), .A2(A[63]), .ZN(n107) );
  OR2_X1 U409 ( .A1(B[60]), .A2(A[60]), .ZN(n129) );
  OR2_X1 U410 ( .A1(A[45]), .A2(B[45]), .ZN(n185) );
  OR2_X1 U411 ( .A1(A[47]), .A2(B[47]), .ZN(n178) );
  AND2_X1 U412 ( .A1(B[34]), .A2(A[34]), .ZN(n77) );
  OR2_X1 U413 ( .A1(B[34]), .A2(A[34]), .ZN(n286) );
  OR2_X1 U414 ( .A1(B[13]), .A2(A[13]), .ZN(n441) );
  INV_X1 U415 ( .A(B[35]), .ZN(n607) );
  INV_X1 U416 ( .A(B[26]), .ZN(n609) );
  INV_X1 U417 ( .A(B[31]), .ZN(n608) );
  OR2_X1 U418 ( .A1(B[6]), .A2(A[6]), .ZN(n98) );
  OR2_X1 U419 ( .A1(B[5]), .A2(A[5]), .ZN(n103) );
  OR2_X1 U420 ( .A1(B[10]), .A2(A[10]), .ZN(n468) );
  OR2_X1 U421 ( .A1(B[9]), .A2(A[9]), .ZN(n85) );
  OR2_X1 U422 ( .A1(B[11]), .A2(A[11]), .ZN(n462) );
  OR2_X1 U423 ( .A1(B[7]), .A2(A[7]), .ZN(n93) );
  OR2_X1 U424 ( .A1(B[8]), .A2(A[8]), .ZN(n89) );
  OR2_X1 U425 ( .A1(B[12]), .A2(A[12]), .ZN(n440) );
  OR2_X1 U426 ( .A1(B[1]), .A2(A[1]), .ZN(n346) );
  OR2_X1 U427 ( .A1(B[2]), .A2(A[2]), .ZN(n348) );
  OR2_X1 U428 ( .A1(B[4]), .A2(A[4]), .ZN(n149) );
  OR2_X1 U429 ( .A1(B[3]), .A2(A[3]), .ZN(n255) );
  OR2_X1 U430 ( .A1(B[0]), .A2(A[0]), .ZN(n481) );
  NAND2_X1 U431 ( .A1(B[1]), .A2(A[1]), .ZN(n345) );
  NAND2_X1 U432 ( .A1(B[8]), .A2(A[8]), .ZN(n90) );
  NAND2_X1 U433 ( .A1(B[12]), .A2(A[12]), .ZN(n433) );
  NAND2_X1 U434 ( .A1(B[13]), .A2(A[13]), .ZN(n434) );
  NAND2_X1 U435 ( .A1(B[6]), .A2(A[6]), .ZN(n95) );
  NAND2_X1 U436 ( .A1(B[9]), .A2(A[9]), .ZN(n86) );
  NAND2_X1 U437 ( .A1(B[2]), .A2(A[2]), .ZN(n253) );
  NAND2_X1 U438 ( .A1(B[0]), .A2(A[0]), .ZN(n413) );
  NAND2_X1 U439 ( .A1(B[4]), .A2(A[4]), .ZN(n148) );
  NAND2_X1 U440 ( .A1(B[5]), .A2(A[5]), .ZN(n102) );
  NAND2_X1 U441 ( .A1(B[10]), .A2(A[10]), .ZN(n465) );
  NAND2_X1 U442 ( .A1(B[3]), .A2(A[3]), .ZN(n256) );
  NAND2_X1 U443 ( .A1(B[7]), .A2(A[7]), .ZN(n94) );
  NAND2_X1 U444 ( .A1(B[11]), .A2(A[11]), .ZN(n466) );
  OR2_X1 U445 ( .A1(B[55]), .A2(A[55]), .ZN(net491458) );
  AND2_X1 U446 ( .A1(B[55]), .A2(A[55]), .ZN(n41) );
  NAND2_X1 U447 ( .A1(A[25]), .A2(B[25]), .ZN(n363) );
  AND2_X1 U448 ( .A1(A[31]), .A2(B[31]), .ZN(n76) );
  NOR2_X1 U449 ( .A1(A[31]), .A2(B[31]), .ZN(n45) );
  OR2_X1 U450 ( .A1(A[31]), .A2(B[31]), .ZN(n44) );
  INV_X1 U451 ( .A(A[31]), .ZN(n579) );
  OAI21_X1 U452 ( .B1(n356), .B2(n357), .A(n61), .ZN(n308) );
  XNOR2_X1 U453 ( .A(n420), .B(n421), .ZN(SUM[17]) );
  XNOR2_X1 U454 ( .A(n210), .B(n209), .ZN(SUM[44]) );
  XNOR2_X1 U455 ( .A(n196), .B(n197), .ZN(SUM[47]) );
  OAI21_X1 U456 ( .B1(n54), .B2(n584), .A(n363), .ZN(n374) );
  INV_X1 U457 ( .A(A[23]), .ZN(n590) );
  NAND2_X1 U458 ( .A1(B[23]), .A2(A[23]), .ZN(n380) );
  INV_X1 U459 ( .A(n143), .ZN(n554) );
  NAND2_X1 U460 ( .A1(n137), .A2(n143), .ZN(n159) );
  NAND2_X1 U461 ( .A1(n239), .A2(n505), .ZN(n233) );
  INV_X1 U462 ( .A(n165), .ZN(n541) );
  NAND2_X1 U463 ( .A1(n165), .A2(n207), .ZN(n210) );
  OR2_X1 U464 ( .A1(net491479), .A2(n531), .ZN(net538270) );
  XNOR2_X1 U465 ( .A(n65), .B(n225), .ZN(SUM[42]) );
  OAI21_X1 U466 ( .B1(n533), .B2(n543), .A(n214), .ZN(n65) );
  OR2_X1 U467 ( .A1(B[27]), .A2(A[27]), .ZN(n61) );
  NAND2_X1 U468 ( .A1(A[27]), .A2(B[27]), .ZN(n360) );
  OR2_X1 U469 ( .A1(A[27]), .A2(B[27]), .ZN(n358) );
  XNOR2_X1 U470 ( .A(net491478), .B(net491475), .ZN(SUM[52]) );
  XNOR2_X1 U471 ( .A(n128), .B(n127), .ZN(SUM[61]) );
  OAI21_X1 U472 ( .B1(n554), .B2(n529), .A(n137), .ZN(n523) );
  INV_X1 U473 ( .A(n246), .ZN(n539) );
  AND2_X1 U474 ( .A1(n246), .A2(n247), .ZN(n239) );
  INV_X1 U475 ( .A(net491492), .ZN(n569) );
  OR2_X1 U476 ( .A1(A[48]), .A2(B[48]), .ZN(net491492) );
  OAI21_X1 U477 ( .B1(n554), .B2(n529), .A(n137), .ZN(n156) );
  NAND4_X1 U478 ( .A1(net491456), .A2(net491457), .A3(net491455), .A4(
        net491458), .ZN(n37) );
  INV_X1 U479 ( .A(net491457), .ZN(n568) );
  NAND2_X1 U480 ( .A1(net491451), .A2(net491457), .ZN(net491473) );
  NAND2_X1 U481 ( .A1(n208), .A2(n195), .ZN(n165) );
  NAND2_X1 U482 ( .A1(n211), .A2(n212), .ZN(n208) );
  NAND2_X1 U483 ( .A1(B[18]), .A2(A[18]), .ZN(n410) );
  NAND2_X1 U484 ( .A1(B[18]), .A2(A[18]), .ZN(n416) );
  AOI21_X1 U485 ( .B1(n1), .B2(n248), .A(n270), .ZN(n267) );
  XNOR2_X1 U486 ( .A(n285), .B(n66), .ZN(SUM[35]) );
  XNOR2_X1 U487 ( .A(net538738), .B(net491504), .ZN(SUM[50]) );
  AND2_X1 U488 ( .A1(n216), .A2(n195), .ZN(n58) );
  AND2_X1 U489 ( .A1(n216), .A2(n217), .ZN(n211) );
  OAI21_X1 U490 ( .B1(n526), .B2(n561), .A(n115), .ZN(n122) );
  INV_X1 U491 ( .A(n127), .ZN(n526) );
  AOI21_X1 U492 ( .B1(n498), .B2(n333), .A(n580), .ZN(n338) );
  NAND2_X1 U493 ( .A1(B[29]), .A2(A[29]), .ZN(n301) );
  OR2_X1 U494 ( .A1(B[29]), .A2(A[29]), .ZN(n81) );
  AOI21_X1 U495 ( .B1(n297), .B2(n298), .A(n76), .ZN(n296) );
  XNOR2_X1 U496 ( .A(net538534), .B(net491511), .ZN(SUM[49]) );
  INV_X1 U497 ( .A(n503), .ZN(n547) );
  AND3_X1 U498 ( .A1(n503), .A2(n177), .A3(n10), .ZN(n72) );
  NAND2_X1 U499 ( .A1(n178), .A2(n177), .ZN(n175) );
  AOI21_X1 U500 ( .B1(n260), .B2(n242), .A(n535), .ZN(n257) );
  NAND2_X1 U501 ( .A1(n242), .A2(n247), .ZN(n262) );
  AND3_X1 U502 ( .A1(n238), .A2(n242), .A3(n19), .ZN(n42) );
  AOI21_X1 U503 ( .B1(n17), .B2(n286), .A(n77), .ZN(n285) );
  AOI21_X1 U504 ( .B1(net491502), .B2(net491491), .A(n571), .ZN(net491497) );
  NAND2_X1 U505 ( .A1(n177), .A2(n183), .ZN(n202) );
  OAI211_X1 U506 ( .C1(n546), .C2(n181), .A(n182), .B(n183), .ZN(n179) );
  AND2_X1 U507 ( .A1(n495), .A2(n192), .ZN(n232) );
  XNOR2_X1 U508 ( .A(n54), .B(n376), .ZN(SUM[25]) );
  OAI21_X1 U509 ( .B1(n525), .B2(n565), .A(net491487), .ZN(net538738) );
  OAI21_X1 U510 ( .B1(n525), .B2(n565), .A(net491487), .ZN(net491502) );
  OAI211_X1 U511 ( .C1(n565), .C2(net491486), .A(net491487), .B(net491488), 
        .ZN(net491483) );
  NAND2_X1 U512 ( .A1(net491487), .A2(net491493), .ZN(net491511) );
  OR2_X1 U513 ( .A1(n16), .A2(n236), .ZN(n14) );
  XNOR2_X1 U514 ( .A(n16), .B(n275), .ZN(SUM[36]) );
  NOR2_X1 U515 ( .A1(n516), .A2(n75), .ZN(n151) );
  NOR2_X1 U516 ( .A1(n556), .A2(n516), .ZN(n134) );
  NAND2_X1 U517 ( .A1(B[60]), .A2(A[60]), .ZN(n116) );
  XNOR2_X1 U518 ( .A(n514), .B(n228), .ZN(SUM[41]) );
  INV_X1 U519 ( .A(n227), .ZN(n533) );
  INV_X1 U520 ( .A(n35), .ZN(n532) );
  OR2_X1 U521 ( .A1(B[59]), .A2(A[59]), .ZN(n145) );
  NAND4_X1 U523 ( .A1(n143), .A2(n144), .A3(n142), .A4(n145), .ZN(n132) );
  NAND2_X1 U525 ( .A1(n67), .A2(n68), .ZN(n340) );
  XNOR2_X1 U526 ( .A(n260), .B(n262), .ZN(SUM[38]) );
  OAI21_X1 U527 ( .B1(n229), .B2(n263), .A(n264), .ZN(n260) );
  XNOR2_X1 U528 ( .A(n523), .B(n157), .ZN(SUM[57]) );
  NOR2_X1 U529 ( .A1(n511), .A2(n566), .ZN(n40) );
  NAND2_X1 U530 ( .A1(n359), .A2(n360), .ZN(n357) );
  AOI211_X1 U531 ( .C1(n609), .C2(n586), .A(n584), .B(n73), .ZN(n356) );
  NAND2_X1 U532 ( .A1(B[56]), .A2(A[56]), .ZN(n137) );
  XNOR2_X1 U534 ( .A(n131), .B(n130), .ZN(SUM[60]) );
  INV_X1 U535 ( .A(n130), .ZN(n527) );
  INV_X1 U536 ( .A(n179), .ZN(n545) );
  OAI21_X1 U537 ( .B1(n132), .B2(n529), .A(n133), .ZN(n130) );
  NAND2_X1 U538 ( .A1(n579), .A2(n608), .ZN(n321) );
  NAND2_X1 U539 ( .A1(n351), .A2(n79), .ZN(n67) );
  AND2_X1 U540 ( .A1(A[51]), .A2(B[51]), .ZN(net534682) );
  OR2_X1 U541 ( .A1(A[51]), .A2(B[51]), .ZN(net491494) );
  OAI21_X1 U542 ( .B1(net491480), .B2(n569), .A(net491486), .ZN(net538534) );
  OAI21_X1 U543 ( .B1(net491480), .B2(n569), .A(net491486), .ZN(net491508) );
  XNOR2_X1 U544 ( .A(net491439), .B(n159), .ZN(SUM[56]) );
  INV_X1 U546 ( .A(net491439), .ZN(n529) );
  NAND2_X1 U547 ( .A1(n512), .A2(n171), .ZN(n169) );
  OAI21_X1 U548 ( .B1(n553), .B2(n170), .A(n272), .ZN(n270) );
  NAND2_X1 U549 ( .A1(A[35]), .A2(B[35]), .ZN(n171) );
  INV_X1 U550 ( .A(A[35]), .ZN(n572) );
  OAI21_X1 U551 ( .B1(n230), .B2(n16), .A(n231), .ZN(n227) );
  NAND2_X1 U552 ( .A1(n42), .A2(n192), .ZN(n230) );
  AOI21_X1 U553 ( .B1(n232), .B2(n64), .A(n550), .ZN(n231) );
  INV_X1 U558 ( .A(n187), .ZN(n524) );
  NOR2_X1 U559 ( .A1(n45), .A2(n581), .ZN(n297) );
  AOI21_X1 U560 ( .B1(n134), .B2(n135), .A(n75), .ZN(n133) );
  NAND2_X1 U561 ( .A1(n418), .A2(n326), .ZN(n417) );
  OAI21_X1 U562 ( .B1(n425), .B2(n426), .A(n427), .ZN(n337) );
  NAND2_X1 U563 ( .A1(B[15]), .A2(A[15]), .ZN(n431) );
  INV_X1 U564 ( .A(net491494), .ZN(n570) );
  AND2_X1 U565 ( .A1(net491494), .A2(net491491), .ZN(net491482) );
  NAND4_X1 U566 ( .A1(net491492), .A2(net491493), .A3(net491491), .A4(
        net491494), .ZN(net491479) );
  OAI211_X1 U567 ( .C1(n49), .C2(n354), .A(n355), .B(n308), .ZN(n9) );
  OAI211_X1 U568 ( .C1(n49), .C2(n354), .A(n355), .B(n308), .ZN(n351) );
  NAND2_X1 U571 ( .A1(n388), .A2(n354), .ZN(n387) );
  OAI21_X1 U572 ( .B1(n26), .B2(n574), .A(n282), .ZN(n17) );
  NAND2_X1 U573 ( .A1(B[48]), .A2(A[48]), .ZN(net491486) );
  NAND2_X1 U575 ( .A1(n9), .A2(n305), .ZN(n342) );
  NAND2_X1 U576 ( .A1(n501), .A2(n359), .ZN(n373) );
  AND4_X1 U577 ( .A1(n358), .A2(n361), .A3(n365), .A4(n501), .ZN(n50) );
  NAND4_X1 U578 ( .A1(n358), .A2(n361), .A3(n365), .A4(n501), .ZN(n49) );
  NAND2_X1 U579 ( .A1(n585), .A2(n362), .ZN(n369) );
  NAND4_X1 U581 ( .A1(n358), .A2(n361), .A3(n365), .A4(n362), .ZN(n353) );
  NAND2_X1 U582 ( .A1(A[43]), .A2(B[43]), .ZN(n216) );
  XNOR2_X1 U583 ( .A(net491497), .B(net491498), .ZN(SUM[51]) );
  NAND2_X1 U584 ( .A1(n161), .A2(n162), .ZN(net491513) );
  AND2_X1 U587 ( .A1(n161), .A2(n162), .ZN(net491480) );
  OAI211_X1 U588 ( .C1(n293), .C2(n294), .A(n502), .B(n496), .ZN(n13) );
  NOR2_X1 U589 ( .A1(n511), .A2(n41), .ZN(net491462) );
  AND3_X1 U590 ( .A1(n512), .A2(n171), .A3(n274), .ZN(n229) );
  AND3_X1 U591 ( .A1(n512), .A2(n171), .A3(n274), .ZN(n16) );
  NAND2_X1 U592 ( .A1(B[17]), .A2(A[17]), .ZN(n409) );
  XNOR2_X1 U593 ( .A(net491461), .B(net491462), .ZN(SUM[55]) );
  XNOR2_X1 U594 ( .A(n510), .B(net491468), .ZN(SUM[54]) );
  AOI21_X1 U595 ( .B1(net491455), .B2(n510), .A(n567), .ZN(net491461) );
  XNOR2_X1 U596 ( .A(n150), .B(n151), .ZN(SUM[59]) );
  XNOR2_X1 U597 ( .A(n152), .B(n154), .ZN(SUM[58]) );
  AOI21_X1 U600 ( .B1(n142), .B2(n152), .A(n555), .ZN(n150) );
  AND2_X1 U601 ( .A1(B[59]), .A2(A[59]), .ZN(n75) );
  AOI21_X1 U602 ( .B1(n172), .B2(n72), .A(n173), .ZN(n161) );
  OAI21_X1 U603 ( .B1(n175), .B2(n545), .A(n176), .ZN(n173) );
  OAI21_X1 U604 ( .B1(n37), .B2(n530), .A(net491445), .ZN(net491439) );
  AOI21_X1 U605 ( .B1(n40), .B2(net491447), .A(n41), .ZN(net491445) );
  OAI21_X1 U606 ( .B1(n528), .B2(n557), .A(n138), .ZN(n152) );
  INV_X1 U607 ( .A(n156), .ZN(n528) );
endmodule


module RCA_NBIT64_9 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_9_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_8_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net492633, net492625, net492611, net492610, net492609, net492608,
         net492604, net492601, net492600, net492589, net492586, net492584,
         net492578, net492577, net492572, net492546, net492533, net492530,
         net492527, net492522, net492520, net492514, net537205, net537537,
         net538271, net538546, net492553, net492532, net492526, net492573,
         net492568, net492567, net492566, net492558, net534634, net492571,
         net538272, net537656, net492563, net492561, net492559, net492555,
         net492574, n2, n3, n4, n7, n9, n10, n11, n12, n13, n14, n15, n16, n18,
         n19, n21, n22, n23, n24, n25, n28, n29, n31, n32, n36, n38, n39, n40,
         n41, n42, n43, n44, n47, n48, n50, n51, n52, n55, n58, n59, n60, n62,
         n63, n64, n67, n68, n69, n70, n71, n73, n74, n77, n78, n79, n81, n83,
         n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n110, n111, n112,
         n113, n115, n116, n117, n118, n119, n120, n122, n123, n126, n127,
         n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n141,
         n142, n143, n144, n145, n146, n147, n148, n151, n152, n153, n154,
         n156, n157, n158, n159, n160, n161, n163, n164, n165, n166, n167,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n196, n197, n198, n199, n201, n204, n206, n209,
         n211, n214, n215, n216, n217, n218, n220, n222, n223, n225, n226,
         n227, n228, n229, n231, n234, n235, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n248, n249, n250, n251, n252, n253,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n280, n281, n282, n283, n284, n285, n286, n287, n290, n291, n292,
         n293, n294, n297, n298, n300, n301, n302, n303, n304, n305, n306,
         n307, n310, n311, n312, n313, n315, n316, n317, n319, n320, n321,
         n322, n323, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n337, n339, n340, n341, n343, n344, n347, n348, n349, n350,
         n352, n353, n354, n355, n356, n357, n359, n360, n361, n362, n363,
         n366, n367, n368, n369, n370, n371, n372, n375, n376, n377, n379,
         n380, n381, n383, n384, n385, n386, n387, n388, n389, n394, n395,
         n396, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n413, n414, n415, n416, n418, n419, n420, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n433, n434,
         n435, n436, n437, n438, n439, n441, n442, n443, n445, n447, n449,
         n450, n453, n454, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n489,
         n490, n491, n492, n494, n496, n497, n498, n499, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622;

  OR2_X2 U7 ( .A1(A[34]), .A2(B[34]), .ZN(n171) );
  NAND3_X1 U9 ( .A1(n167), .A2(n169), .A3(n4), .ZN(n157) );
  NAND3_X1 U17 ( .A1(n182), .A2(n73), .A3(n3), .ZN(n22) );
  OR2_X2 U18 ( .A1(B[46]), .A2(A[46]), .ZN(n169) );
  XOR2_X1 U46 ( .A(n24), .B(n426), .Z(SUM[19]) );
  NAND3_X1 U62 ( .A1(n619), .A2(n547), .A3(n307), .ZN(n359) );
  NAND3_X1 U72 ( .A1(n566), .A2(n277), .A3(n69), .ZN(n271) );
  NAND3_X1 U75 ( .A1(n235), .A2(n238), .A3(n518), .ZN(n237) );
  OR2_X2 U76 ( .A1(A[44]), .A2(B[44]), .ZN(n172) );
  NAND3_X1 U81 ( .A1(n238), .A2(n518), .A3(n235), .ZN(n231) );
  NAND3_X1 U84 ( .A1(n353), .A2(n355), .A3(n354), .ZN(n340) );
  XOR2_X1 U185 ( .A(n218), .B(n83), .Z(SUM[44]) );
  OR2_X2 U374 ( .A1(A[29]), .A2(B[29]), .ZN(n320) );
  OR2_X2 U394 ( .A1(B[36]), .A2(A[36]), .ZN(n253) );
  NAND3_X1 U549 ( .A1(n190), .A2(n10), .A3(n192), .ZN(n189) );
  NAND3_X1 U560 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n238) );
  NAND3_X1 U563 ( .A1(n198), .A2(n271), .A3(n272), .ZN(n270) );
  NAND3_X1 U570 ( .A1(n173), .A2(n179), .A3(n178), .ZN(n291) );
  NAND3_X1 U584 ( .A1(n319), .A2(n360), .A3(n18), .ZN(n353) );
  NAND3_X1 U589 ( .A1(n305), .A2(n306), .A3(n307), .ZN(n356) );
  NAND3_X1 U594 ( .A1(n385), .A2(n370), .A3(n384), .ZN(n379) );
  NAND3_X1 U595 ( .A1(n327), .A2(n64), .A3(n404), .ZN(n395) );
  NAND3_X1 U619 ( .A1(n477), .A2(n478), .A3(n479), .ZN(n476) );
  NAND3_X1 U620 ( .A1(n480), .A2(n93), .A3(n481), .ZN(n477) );
  OR2_X2 U120 ( .A1(B[54]), .A2(A[54]), .ZN(net492571) );
  OR2_X2 U132 ( .A1(B[56]), .A2(A[56]), .ZN(n52) );
  OR2_X2 U141 ( .A1(B[57]), .A2(A[57]), .ZN(net492532) );
  OR2_X2 U189 ( .A1(B[45]), .A2(A[45]), .ZN(n174) );
  OR2_X2 U387 ( .A1(B[32]), .A2(A[32]), .ZN(n179) );
  OR2_X2 U391 ( .A1(B[58]), .A2(A[58]), .ZN(net492530) );
  OR2_X2 U402 ( .A1(B[48]), .A2(A[48]), .ZN(net492604) );
  OR2_X2 U418 ( .A1(B[50]), .A2(A[50]), .ZN(net492600) );
  AND2_X1 U2 ( .A1(n327), .A2(n403), .ZN(n389) );
  INV_X1 U3 ( .A(n164), .ZN(n591) );
  OR2_X1 U4 ( .A1(A[49]), .A2(B[49]), .ZN(net492625) );
  OR2_X1 U5 ( .A1(A[51]), .A2(B[51]), .ZN(net492601) );
  AND2_X1 U6 ( .A1(n494), .A2(n425), .ZN(SUM[0]) );
  OR2_X1 U8 ( .A1(A[59]), .A2(B[59]), .ZN(net492533) );
  CLKBUF_X1 U10 ( .A(A[24]), .Z(n502) );
  AND2_X1 U11 ( .A1(net492573), .A2(net492572), .ZN(n503) );
  XNOR2_X1 U12 ( .A(n533), .B(n504), .ZN(SUM[42]) );
  AND2_X1 U13 ( .A1(n523), .A2(n186), .ZN(n504) );
  OR2_X1 U14 ( .A1(A[38]), .A2(B[38]), .ZN(n252) );
  OAI21_X1 U15 ( .B1(n541), .B2(n581), .A(net492526), .ZN(n505) );
  XNOR2_X1 U16 ( .A(n506), .B(n507), .ZN(SUM[33]) );
  AND2_X1 U19 ( .A1(n297), .A2(n283), .ZN(n506) );
  AND2_X1 U20 ( .A1(n284), .A2(n178), .ZN(n507) );
  CLKBUF_X1 U21 ( .A(n307), .Z(n508) );
  AND2_X1 U22 ( .A1(n271), .A2(n199), .ZN(n509) );
  CLKBUF_X1 U23 ( .A(net492567), .Z(n510) );
  AND2_X1 U24 ( .A1(n271), .A2(n199), .ZN(n511) );
  AND2_X1 U25 ( .A1(n42), .A2(n43), .ZN(n512) );
  AND2_X1 U26 ( .A1(n42), .A2(n43), .ZN(net537656) );
  CLKBUF_X1 U27 ( .A(n306), .Z(n513) );
  AND2_X1 U28 ( .A1(n368), .A2(n372), .ZN(n514) );
  AND3_X1 U29 ( .A1(n366), .A2(n371), .A3(n514), .ZN(n18) );
  OR2_X2 U30 ( .A1(A[25]), .A2(B[25]), .ZN(n368) );
  OR2_X2 U31 ( .A1(A[22]), .A2(B[22]), .ZN(n327) );
  NAND3_X1 U32 ( .A1(net492574), .A2(net492571), .A3(n503), .ZN(net492559) );
  NOR2_X1 U33 ( .A1(B[55]), .A2(A[55]), .ZN(n515) );
  OR2_X1 U34 ( .A1(B[52]), .A2(A[52]), .ZN(net492572) );
  OR2_X1 U35 ( .A1(A[53]), .A2(B[53]), .ZN(net492573) );
  OR2_X1 U36 ( .A1(B[39]), .A2(A[39]), .ZN(n10) );
  NAND2_X1 U37 ( .A1(n291), .A2(n290), .ZN(n516) );
  OR2_X1 U38 ( .A1(n62), .A2(n177), .ZN(n517) );
  OR2_X2 U39 ( .A1(A[33]), .A2(B[33]), .ZN(n178) );
  BUF_X1 U40 ( .A(n222), .Z(n518) );
  NAND3_X1 U41 ( .A1(n353), .A2(n355), .A3(n354), .ZN(n519) );
  OR2_X1 U42 ( .A1(n40), .A2(n175), .ZN(n520) );
  OR2_X1 U43 ( .A1(n40), .A2(n175), .ZN(n225) );
  OR2_X1 U44 ( .A1(A[43]), .A2(B[43]), .ZN(n521) );
  OR2_X1 U45 ( .A1(A[43]), .A2(B[43]), .ZN(n187) );
  AND2_X1 U47 ( .A1(net492574), .A2(net492571), .ZN(n41) );
  NAND2_X1 U48 ( .A1(n265), .A2(n266), .ZN(n522) );
  CLKBUF_X1 U49 ( .A(n31), .Z(n523) );
  OR2_X1 U50 ( .A1(A[42]), .A2(B[42]), .ZN(n186) );
  OR2_X1 U51 ( .A1(n222), .A2(n28), .ZN(n524) );
  NAND2_X1 U52 ( .A1(n525), .A2(n524), .ZN(n29) );
  AND2_X1 U53 ( .A1(n31), .A2(n223), .ZN(n525) );
  AND2_X1 U54 ( .A1(net538272), .A2(net492561), .ZN(n526) );
  XNOR2_X1 U55 ( .A(n522), .B(n527), .ZN(SUM[38]) );
  NAND2_X1 U56 ( .A1(n252), .A2(n264), .ZN(n527) );
  XNOR2_X1 U57 ( .A(n201), .B(n528), .ZN(SUM[47]) );
  NOR2_X1 U58 ( .A1(n87), .A2(n590), .ZN(n528) );
  XOR2_X1 U59 ( .A(n237), .B(n529), .Z(SUM[41]) );
  AND2_X1 U60 ( .A1(n223), .A2(n597), .ZN(n529) );
  XOR2_X1 U61 ( .A(n530), .B(n535), .Z(SUM[50]) );
  NAND2_X1 U63 ( .A1(net492600), .A2(net492611), .ZN(n530) );
  XOR2_X1 U64 ( .A(n512), .B(n531), .Z(SUM[52]) );
  NAND2_X1 U65 ( .A1(net492572), .A2(net492566), .ZN(n531) );
  XOR2_X1 U66 ( .A(net537537), .B(n532), .Z(SUM[48]) );
  AND2_X1 U67 ( .A1(net492604), .A2(net492609), .ZN(n532) );
  AND2_X1 U68 ( .A1(n234), .A2(n223), .ZN(n533) );
  INV_X1 U69 ( .A(n403), .ZN(n561) );
  XNOR2_X1 U70 ( .A(n19), .B(n383), .ZN(SUM[25]) );
  NOR2_X1 U71 ( .A1(n550), .A2(n549), .ZN(n383) );
  NOR2_X1 U73 ( .A1(n594), .A2(n29), .ZN(n183) );
  NAND2_X1 U74 ( .A1(n520), .A2(n226), .ZN(n243) );
  INV_X1 U77 ( .A(A[27]), .ZN(n552) );
  INV_X1 U78 ( .A(n177), .ZN(n592) );
  INV_X1 U79 ( .A(n316), .ZN(n544) );
  AND2_X1 U80 ( .A1(n356), .A2(n310), .ZN(n16) );
  OAI21_X1 U82 ( .B1(n620), .B2(n461), .A(n458), .ZN(n96) );
  AOI21_X1 U83 ( .B1(n457), .B2(n458), .A(n459), .ZN(n454) );
  NAND2_X1 U85 ( .A1(n614), .A2(n460), .ZN(n457) );
  INV_X1 U86 ( .A(n461), .ZN(n614) );
  NAND4_X1 U87 ( .A1(n89), .A2(n563), .A3(n18), .A4(n317), .ZN(n301) );
  INV_X1 U88 ( .A(n323), .ZN(n563) );
  NOR2_X1 U89 ( .A1(n603), .A2(n316), .ZN(n317) );
  NAND2_X1 U90 ( .A1(n474), .A2(n456), .ZN(n472) );
  NAND2_X1 U91 ( .A1(n610), .A2(n96), .ZN(n474) );
  INV_X1 U92 ( .A(n459), .ZN(n610) );
  INV_X1 U93 ( .A(n423), .ZN(n603) );
  INV_X1 U94 ( .A(n460), .ZN(n620) );
  NOR2_X1 U95 ( .A1(n113), .A2(n576), .ZN(SUM[64]) );
  INV_X1 U96 ( .A(n456), .ZN(n611) );
  NOR2_X1 U97 ( .A1(n560), .A2(n559), .ZN(n344) );
  INV_X1 U98 ( .A(n332), .ZN(n560) );
  XNOR2_X1 U99 ( .A(n337), .B(n60), .ZN(SUM[31]) );
  NOR2_X1 U100 ( .A1(n558), .A2(n557), .ZN(n60) );
  AOI21_X1 U101 ( .B1(n339), .B2(n519), .A(n341), .ZN(n337) );
  INV_X1 U102 ( .A(n331), .ZN(n558) );
  OR2_X1 U103 ( .A1(n587), .A2(n588), .ZN(n83) );
  AOI21_X1 U104 ( .B1(n592), .B2(n243), .A(n220), .ZN(n218) );
  AND2_X1 U105 ( .A1(n169), .A2(n12), .ZN(n3) );
  NAND2_X1 U106 ( .A1(n388), .A2(n327), .ZN(n409) );
  NAND2_X1 U107 ( .A1(n52), .A2(n51), .ZN(net492558) );
  NAND2_X1 U108 ( .A1(n310), .A2(n508), .ZN(n32) );
  OAI21_X1 U109 ( .B1(n376), .B2(n377), .A(n513), .ZN(n375) );
  NAND2_X1 U110 ( .A1(n368), .A2(n63), .ZN(n377) );
  INV_X1 U111 ( .A(net492527), .ZN(n579) );
  NAND2_X1 U112 ( .A1(n399), .A2(n328), .ZN(n405) );
  NAND4_X1 U113 ( .A1(net492533), .A2(net492532), .A3(net492530), .A4(n52), 
        .ZN(n50) );
  AOI21_X1 U114 ( .B1(n416), .B2(n427), .A(n600), .ZN(n426) );
  NAND2_X1 U115 ( .A1(n422), .A2(n414), .ZN(n24) );
  OAI21_X1 U116 ( .B1(n71), .B2(n571), .A(net492611), .ZN(n148) );
  INV_X1 U117 ( .A(net492568), .ZN(n583) );
  XNOR2_X1 U118 ( .A(n381), .B(n380), .ZN(SUM[26]) );
  NAND2_X1 U119 ( .A1(n63), .A2(n306), .ZN(n380) );
  OAI21_X1 U121 ( .B1(n19), .B2(n550), .A(n369), .ZN(n381) );
  AND2_X1 U122 ( .A1(n319), .A2(n359), .ZN(n357) );
  XNOR2_X1 U123 ( .A(n64), .B(n411), .ZN(SUM[20]) );
  NAND2_X1 U124 ( .A1(n325), .A2(n402), .ZN(n411) );
  INV_X1 U125 ( .A(n21), .ZN(n539) );
  NAND2_X1 U126 ( .A1(net492571), .A2(net492568), .ZN(net492584) );
  NAND2_X1 U127 ( .A1(net492530), .A2(net492527), .ZN(n145) );
  XNOR2_X1 U128 ( .A(n242), .B(n243), .ZN(SUM[40]) );
  XOR2_X1 U129 ( .A(n40), .B(n276), .Z(SUM[36]) );
  AOI21_X1 U130 ( .B1(n311), .B2(n312), .A(n313), .ZN(n303) );
  AND2_X1 U131 ( .A1(n304), .A2(n356), .ZN(n13) );
  XNOR2_X1 U133 ( .A(n516), .B(n292), .ZN(SUM[34]) );
  NAND2_X1 U134 ( .A1(n171), .A2(n285), .ZN(n292) );
  OAI21_X1 U135 ( .B1(n386), .B2(n396), .A(n387), .ZN(n311) );
  XNOR2_X1 U136 ( .A(n154), .B(net492633), .ZN(SUM[49]) );
  NOR2_X1 U137 ( .A1(n572), .A2(n573), .ZN(net492633) );
  NAND2_X1 U138 ( .A1(n367), .A2(n368), .ZN(n305) );
  NAND2_X1 U139 ( .A1(n369), .A2(n370), .ZN(n367) );
  XNOR2_X1 U140 ( .A(n340), .B(n352), .ZN(SUM[29]) );
  NAND2_X1 U142 ( .A1(n320), .A2(n334), .ZN(n352) );
  NAND2_X1 U143 ( .A1(n331), .A2(n332), .ZN(n330) );
  AOI21_X1 U144 ( .B1(n333), .B2(n334), .A(n559), .ZN(n329) );
  NAND2_X1 U145 ( .A1(n553), .A2(n320), .ZN(n333) );
  XNOR2_X1 U146 ( .A(n298), .B(n69), .ZN(SUM[32]) );
  NAND2_X1 U147 ( .A1(n179), .A2(n283), .ZN(n298) );
  XNOR2_X1 U148 ( .A(n55), .B(n410), .ZN(SUM[21]) );
  NAND2_X1 U149 ( .A1(n326), .A2(n401), .ZN(n410) );
  OAI21_X1 U150 ( .B1(n561), .B2(n546), .A(n402), .ZN(n55) );
  INV_X1 U151 ( .A(n325), .ZN(n546) );
  XNOR2_X1 U152 ( .A(n361), .B(n362), .ZN(SUM[28]) );
  NOR2_X1 U153 ( .A1(n553), .A2(n554), .ZN(n362) );
  AOI21_X1 U154 ( .B1(n18), .B2(n360), .A(n363), .ZN(n361) );
  INV_X1 U155 ( .A(n319), .ZN(n554) );
  NAND4_X1 U156 ( .A1(n325), .A2(n326), .A3(n327), .A4(n328), .ZN(n316) );
  XNOR2_X1 U157 ( .A(n286), .B(n287), .ZN(SUM[35]) );
  NOR2_X1 U158 ( .A1(n569), .A2(n70), .ZN(n287) );
  AOI21_X1 U159 ( .B1(n293), .B2(n171), .A(n565), .ZN(n286) );
  INV_X1 U160 ( .A(n199), .ZN(n569) );
  XNOR2_X1 U161 ( .A(n58), .B(n206), .ZN(SUM[46]) );
  NAND2_X1 U162 ( .A1(n169), .A2(n164), .ZN(n206) );
  OAI21_X1 U163 ( .B1(n589), .B2(n7), .A(n165), .ZN(n58) );
  OAI211_X1 U164 ( .C1(n396), .C2(n386), .A(n387), .B(n372), .ZN(n385) );
  OAI211_X1 U165 ( .C1(n573), .C2(net492609), .A(net492610), .B(net492611), 
        .ZN(n48) );
  AOI21_X1 U166 ( .B1(n215), .B2(n216), .A(n595), .ZN(n220) );
  NAND3_X1 U167 ( .A1(n521), .A2(n186), .A3(n2), .ZN(n177) );
  AND2_X1 U168 ( .A1(n597), .A2(n79), .ZN(n2) );
  OAI21_X1 U169 ( .B1(n543), .B2(n38), .A(n401), .ZN(n408) );
  INV_X1 U170 ( .A(n326), .ZN(n543) );
  AOI21_X1 U171 ( .B1(n403), .B2(n325), .A(n545), .ZN(n38) );
  INV_X1 U172 ( .A(n402), .ZN(n545) );
  XNOR2_X1 U173 ( .A(n429), .B(n427), .ZN(SUM[18]) );
  NAND2_X1 U174 ( .A1(n416), .A2(n428), .ZN(n429) );
  NAND2_X1 U175 ( .A1(n618), .A2(n552), .ZN(n310) );
  XNOR2_X1 U176 ( .A(n534), .B(n7), .ZN(SUM[45]) );
  AND2_X1 U177 ( .A1(n165), .A2(n174), .ZN(n534) );
  XNOR2_X1 U178 ( .A(net492589), .B(net537205), .ZN(SUM[53]) );
  OAI21_X1 U179 ( .B1(n584), .B2(n512), .A(net492566), .ZN(net537205) );
  AOI21_X1 U180 ( .B1(n215), .B2(n216), .A(n217), .ZN(n214) );
  INV_X1 U181 ( .A(n321), .ZN(n559) );
  NAND4_X1 U182 ( .A1(n192), .A2(n79), .A3(n10), .A4(n190), .ZN(n235) );
  OAI21_X1 U183 ( .B1(n334), .B2(n559), .A(n332), .ZN(n341) );
  NAND2_X1 U184 ( .A1(n395), .A2(n311), .ZN(n360) );
  AND3_X1 U186 ( .A1(n328), .A2(n326), .A3(n325), .ZN(n404) );
  AOI21_X1 U187 ( .B1(n47), .B2(n48), .A(n570), .ZN(n42) );
  NOR2_X1 U188 ( .A1(n573), .A2(n586), .ZN(n44) );
  AOI21_X1 U190 ( .B1(n548), .B2(n508), .A(n551), .ZN(n304) );
  INV_X1 U191 ( .A(n366), .ZN(n548) );
  INV_X1 U192 ( .A(n310), .ZN(n551) );
  NAND4_X1 U193 ( .A1(n371), .A2(n372), .A3(n368), .A4(n366), .ZN(n313) );
  AND2_X1 U194 ( .A1(n152), .A2(n151), .ZN(n535) );
  AND2_X1 U195 ( .A1(n170), .A2(n564), .ZN(n4) );
  INV_X1 U196 ( .A(n175), .ZN(n564) );
  NOR2_X1 U197 ( .A1(n70), .A2(n567), .ZN(n280) );
  INV_X1 U198 ( .A(n171), .ZN(n567) );
  AND2_X1 U199 ( .A1(n191), .A2(n252), .ZN(n241) );
  NOR2_X1 U200 ( .A1(n77), .A2(n78), .ZN(n239) );
  INV_X1 U201 ( .A(n28), .ZN(n597) );
  AND2_X1 U202 ( .A1(n356), .A2(n536), .ZN(n363) );
  AND2_X1 U203 ( .A1(n359), .A2(n310), .ZN(n536) );
  NOR2_X1 U204 ( .A1(n556), .A2(n559), .ZN(n339) );
  INV_X1 U205 ( .A(n320), .ZN(n556) );
  NOR2_X1 U206 ( .A1(n549), .A2(n379), .ZN(n376) );
  OAI21_X1 U207 ( .B1(n596), .B2(n223), .A(n523), .ZN(n229) );
  INV_X1 U208 ( .A(net492625), .ZN(n573) );
  AND3_X1 U209 ( .A1(n385), .A2(n370), .A3(n384), .ZN(n19) );
  NAND2_X1 U210 ( .A1(n291), .A2(n290), .ZN(n293) );
  NAND2_X1 U211 ( .A1(n294), .A2(n178), .ZN(n290) );
  AND3_X1 U212 ( .A1(n327), .A2(n400), .A3(n326), .ZN(n386) );
  NAND2_X1 U213 ( .A1(n401), .A2(n402), .ZN(n400) );
  NAND2_X1 U214 ( .A1(n399), .A2(n388), .ZN(n396) );
  INV_X1 U215 ( .A(n174), .ZN(n589) );
  NAND2_X1 U216 ( .A1(n265), .A2(n266), .ZN(n268) );
  NAND2_X1 U217 ( .A1(n270), .A2(n269), .ZN(n265) );
  NOR2_X1 U218 ( .A1(n9), .A2(n593), .ZN(n269) );
  NAND2_X1 U219 ( .A1(n552), .A2(n618), .ZN(n371) );
  NAND2_X1 U220 ( .A1(n231), .A2(n597), .ZN(n234) );
  XNOR2_X1 U221 ( .A(n274), .B(n273), .ZN(SUM[37]) );
  NAND2_X1 U222 ( .A1(n266), .A2(n197), .ZN(n273) );
  NAND2_X1 U223 ( .A1(n275), .A2(n249), .ZN(n274) );
  AND3_X1 U224 ( .A1(n322), .A2(n320), .A3(n59), .ZN(n89) );
  AND2_X1 U225 ( .A1(n321), .A2(n319), .ZN(n59) );
  INV_X1 U226 ( .A(n216), .ZN(n594) );
  OAI21_X1 U227 ( .B1(n584), .B2(net537656), .A(net492566), .ZN(net492586) );
  INV_X1 U228 ( .A(n368), .ZN(n550) );
  INV_X1 U229 ( .A(n369), .ZN(n549) );
  INV_X1 U230 ( .A(n322), .ZN(n557) );
  AND2_X1 U231 ( .A1(n433), .A2(n418), .ZN(n430) );
  NAND2_X1 U232 ( .A1(n423), .A2(n420), .ZN(n433) );
  INV_X1 U233 ( .A(n354), .ZN(n553) );
  INV_X1 U234 ( .A(n428), .ZN(n600) );
  NAND2_X1 U235 ( .A1(n193), .A2(n194), .ZN(n188) );
  NOR2_X1 U236 ( .A1(n593), .A2(n196), .ZN(n194) );
  NAND2_X1 U237 ( .A1(n191), .A2(n197), .ZN(n196) );
  INV_X1 U238 ( .A(net492572), .ZN(n584) );
  INV_X1 U239 ( .A(n252), .ZN(n599) );
  INV_X1 U240 ( .A(n136), .ZN(n578) );
  INV_X1 U241 ( .A(net492573), .ZN(n574) );
  OR2_X1 U242 ( .A1(n36), .A2(n537), .ZN(n384) );
  NAND2_X1 U243 ( .A1(n389), .A2(n328), .ZN(n537) );
  OR2_X1 U244 ( .A1(n180), .A2(n181), .ZN(n73) );
  AOI21_X1 U245 ( .B1(n188), .B2(n189), .A(n177), .ZN(n180) );
  NOR2_X1 U246 ( .A1(n183), .A2(n184), .ZN(n181) );
  INV_X1 U247 ( .A(n187), .ZN(n595) );
  INV_X1 U248 ( .A(n133), .ZN(n577) );
  INV_X1 U249 ( .A(n129), .ZN(n575) );
  INV_X1 U250 ( .A(n163), .ZN(n587) );
  INV_X1 U251 ( .A(n158), .ZN(n590) );
  NAND2_X1 U252 ( .A1(n146), .A2(n25), .ZN(n152) );
  NAND4_X1 U253 ( .A1(n157), .A2(n156), .A3(n158), .A4(n159), .ZN(n146) );
  AND2_X1 U254 ( .A1(net492625), .A2(net492604), .ZN(n25) );
  NAND4_X1 U255 ( .A1(n182), .A2(n169), .A3(n73), .A4(n12), .ZN(n156) );
  INV_X1 U256 ( .A(net492609), .ZN(n585) );
  INV_X1 U257 ( .A(n264), .ZN(n598) );
  INV_X1 U258 ( .A(n52), .ZN(n582) );
  NAND2_X1 U259 ( .A1(n244), .A2(n192), .ZN(n226) );
  AND2_X1 U260 ( .A1(n10), .A2(n11), .ZN(n244) );
  INV_X1 U261 ( .A(net492608), .ZN(n570) );
  NAND2_X1 U262 ( .A1(n225), .A2(n226), .ZN(n211) );
  INV_X1 U263 ( .A(net492532), .ZN(n581) );
  INV_X1 U264 ( .A(net492604), .ZN(n586) );
  INV_X1 U265 ( .A(n285), .ZN(n565) );
  INV_X1 U266 ( .A(n334), .ZN(n555) );
  AND2_X1 U267 ( .A1(n249), .A2(n199), .ZN(n272) );
  AND2_X1 U268 ( .A1(n174), .A2(n88), .ZN(n170) );
  INV_X1 U269 ( .A(n70), .ZN(n568) );
  XNOR2_X1 U270 ( .A(n430), .B(n431), .ZN(SUM[17]) );
  INV_X1 U271 ( .A(n419), .ZN(n602) );
  XNOR2_X1 U272 ( .A(n470), .B(n469), .ZN(SUM[13]) );
  NAND2_X1 U273 ( .A1(n447), .A2(n449), .ZN(n470) );
  XNOR2_X1 U274 ( .A(n462), .B(n463), .ZN(SUM[15]) );
  NAND2_X1 U275 ( .A1(n464), .A2(n443), .ZN(n463) );
  NAND2_X1 U276 ( .A1(n441), .A2(n439), .ZN(n462) );
  NAND2_X1 U277 ( .A1(n445), .A2(n465), .ZN(n464) );
  XNOR2_X1 U278 ( .A(n434), .B(n423), .ZN(SUM[16]) );
  NAND2_X1 U279 ( .A1(n420), .A2(n418), .ZN(n434) );
  XNOR2_X1 U280 ( .A(n466), .B(n465), .ZN(SUM[14]) );
  NAND2_X1 U281 ( .A1(n445), .A2(n443), .ZN(n466) );
  XNOR2_X1 U282 ( .A(n99), .B(n100), .ZN(SUM[7]) );
  NAND2_X1 U283 ( .A1(n103), .A2(n104), .ZN(n99) );
  NAND2_X1 U284 ( .A1(n101), .A2(n102), .ZN(n100) );
  NAND2_X1 U285 ( .A1(n105), .A2(n106), .ZN(n104) );
  XNOR2_X1 U286 ( .A(n255), .B(n256), .ZN(SUM[3]) );
  NAND2_X1 U287 ( .A1(n259), .A2(n260), .ZN(n255) );
  NAND2_X1 U288 ( .A1(n257), .A2(n258), .ZN(n256) );
  NAND2_X1 U289 ( .A1(n261), .A2(n262), .ZN(n260) );
  XNOR2_X1 U290 ( .A(n482), .B(n483), .ZN(SUM[11]) );
  NAND2_X1 U291 ( .A1(n478), .A2(n484), .ZN(n483) );
  NAND2_X1 U292 ( .A1(n479), .A2(n475), .ZN(n482) );
  NAND2_X1 U293 ( .A1(n481), .A2(n485), .ZN(n484) );
  XNOR2_X1 U294 ( .A(n424), .B(n622), .ZN(SUM[1]) );
  NAND2_X1 U295 ( .A1(n350), .A2(n349), .ZN(n424) );
  XNOR2_X1 U296 ( .A(n95), .B(n96), .ZN(SUM[8]) );
  NAND2_X1 U297 ( .A1(n97), .A2(n98), .ZN(n95) );
  XNOR2_X1 U298 ( .A(n473), .B(n472), .ZN(SUM[12]) );
  NAND2_X1 U299 ( .A1(n453), .A2(n450), .ZN(n473) );
  XNOR2_X1 U300 ( .A(n91), .B(n92), .ZN(SUM[9]) );
  NAND2_X1 U301 ( .A1(n93), .A2(n94), .ZN(n91) );
  XNOR2_X1 U302 ( .A(n139), .B(n112), .ZN(SUM[5]) );
  NAND2_X1 U303 ( .A1(n111), .A2(n110), .ZN(n139) );
  XNOR2_X1 U304 ( .A(n107), .B(n105), .ZN(SUM[6]) );
  NAND2_X1 U305 ( .A1(n106), .A2(n103), .ZN(n107) );
  XNOR2_X1 U306 ( .A(n486), .B(n485), .ZN(SUM[10]) );
  NAND2_X1 U307 ( .A1(n481), .A2(n478), .ZN(n486) );
  XNOR2_X1 U308 ( .A(n347), .B(n261), .ZN(SUM[2]) );
  NAND2_X1 U309 ( .A1(n262), .A2(n259), .ZN(n347) );
  XNOR2_X1 U310 ( .A(n153), .B(n460), .ZN(SUM[4]) );
  NAND2_X1 U311 ( .A1(n142), .A2(n141), .ZN(n153) );
  OAI21_X1 U312 ( .B1(n496), .B2(n497), .A(n258), .ZN(n460) );
  NAND2_X1 U313 ( .A1(n262), .A2(n257), .ZN(n497) );
  NOR2_X1 U314 ( .A1(n498), .A2(n499), .ZN(n496) );
  NAND2_X1 U315 ( .A1(n259), .A2(n349), .ZN(n499) );
  OAI21_X1 U316 ( .B1(n435), .B2(n436), .A(n437), .ZN(n423) );
  NOR2_X1 U317 ( .A1(n454), .A2(n611), .ZN(n435) );
  NAND4_X1 U318 ( .A1(n453), .A2(n447), .A3(n445), .A4(n439), .ZN(n436) );
  AOI21_X1 U319 ( .B1(n438), .B2(n439), .A(n604), .ZN(n437) );
  OAI21_X1 U320 ( .B1(n613), .B2(n612), .A(n94), .ZN(n485) );
  INV_X1 U321 ( .A(n92), .ZN(n613) );
  INV_X1 U322 ( .A(n93), .ZN(n612) );
  OAI21_X1 U323 ( .B1(n608), .B2(n606), .A(n449), .ZN(n465) );
  INV_X1 U324 ( .A(n469), .ZN(n608) );
  INV_X1 U325 ( .A(n447), .ZN(n606) );
  OAI21_X1 U326 ( .B1(n617), .B2(n620), .A(n141), .ZN(n112) );
  INV_X1 U327 ( .A(n142), .ZN(n617) );
  OAI21_X1 U328 ( .B1(n616), .B2(n615), .A(n110), .ZN(n105) );
  INV_X1 U329 ( .A(n112), .ZN(n616) );
  INV_X1 U330 ( .A(n111), .ZN(n615) );
  OAI21_X1 U331 ( .B1(n490), .B2(n491), .A(n101), .ZN(n458) );
  NAND2_X1 U332 ( .A1(n102), .A2(n103), .ZN(n491) );
  NOR2_X1 U333 ( .A1(n15), .A2(n492), .ZN(n490) );
  AND2_X1 U334 ( .A1(n110), .A2(n141), .ZN(n15) );
  NAND4_X1 U335 ( .A1(n420), .A2(n601), .A3(n416), .A4(n422), .ZN(n323) );
  NAND4_X1 U336 ( .A1(n142), .A2(n111), .A3(n106), .A4(n101), .ZN(n461) );
  NAND4_X1 U337 ( .A1(n93), .A2(n97), .A3(n481), .A4(n475), .ZN(n459) );
  AOI21_X1 U338 ( .B1(n116), .B2(n117), .A(n118), .ZN(n113) );
  NAND2_X1 U339 ( .A1(n119), .A2(n120), .ZN(n118) );
  NOR2_X1 U340 ( .A1(n575), .A2(n577), .ZN(n116) );
  AOI21_X1 U341 ( .B1(n442), .B2(n443), .A(n605), .ZN(n438) );
  INV_X1 U342 ( .A(n445), .ZN(n605) );
  AOI21_X1 U343 ( .B1(n609), .B2(n447), .A(n607), .ZN(n442) );
  INV_X1 U344 ( .A(n449), .ZN(n607) );
  NOR2_X1 U345 ( .A1(n621), .A2(n425), .ZN(n498) );
  INV_X1 U346 ( .A(n350), .ZN(n621) );
  NAND2_X1 U347 ( .A1(n489), .A2(n98), .ZN(n92) );
  NAND2_X1 U348 ( .A1(n96), .A2(n97), .ZN(n489) );
  NAND2_X1 U349 ( .A1(n471), .A2(n450), .ZN(n469) );
  NAND2_X1 U350 ( .A1(n472), .A2(n453), .ZN(n471) );
  NAND2_X1 U351 ( .A1(n348), .A2(n349), .ZN(n261) );
  NAND2_X1 U352 ( .A1(n350), .A2(n622), .ZN(n348) );
  NAND2_X1 U353 ( .A1(n475), .A2(n476), .ZN(n456) );
  NAND2_X1 U354 ( .A1(n94), .A2(n98), .ZN(n480) );
  INV_X1 U355 ( .A(n425), .ZN(n622) );
  NAND2_X1 U356 ( .A1(n111), .A2(n106), .ZN(n492) );
  INV_X1 U357 ( .A(n450), .ZN(n609) );
  INV_X1 U358 ( .A(n441), .ZN(n604) );
  NOR2_X1 U359 ( .A1(B[35]), .A2(A[35]), .ZN(n70) );
  NOR2_X1 U360 ( .A1(A[19]), .A2(B[19]), .ZN(n67) );
  AOI21_X1 U361 ( .B1(n416), .B2(n415), .A(n600), .ZN(n413) );
  OR2_X1 U362 ( .A1(A[20]), .A2(B[20]), .ZN(n325) );
  OR2_X1 U363 ( .A1(A[21]), .A2(B[21]), .ZN(n326) );
  NAND2_X1 U364 ( .A1(A[20]), .A2(B[20]), .ZN(n402) );
  NAND2_X1 U365 ( .A1(B[41]), .A2(A[41]), .ZN(n223) );
  NAND2_X1 U366 ( .A1(B[29]), .A2(A[29]), .ZN(n334) );
  NOR2_X1 U367 ( .A1(B[41]), .A2(A[41]), .ZN(n28) );
  NAND2_X1 U368 ( .A1(A[24]), .A2(B[24]), .ZN(n370) );
  XNOR2_X1 U369 ( .A(n394), .B(n360), .ZN(SUM[24]) );
  NAND2_X1 U370 ( .A1(n14), .A2(n370), .ZN(n394) );
  OR2_X1 U371 ( .A1(B[24]), .A2(n502), .ZN(n14) );
  NAND2_X1 U372 ( .A1(A[27]), .A2(B[27]), .ZN(n307) );
  INV_X1 U373 ( .A(B[26]), .ZN(n619) );
  INV_X1 U375 ( .A(A[26]), .ZN(n547) );
  NAND2_X1 U376 ( .A1(B[45]), .A2(A[45]), .ZN(n165) );
  OR2_X1 U377 ( .A1(A[18]), .A2(B[18]), .ZN(n416) );
  AND2_X1 U378 ( .A1(n178), .A2(n179), .ZN(n277) );
  INV_X1 U379 ( .A(n39), .ZN(n566) );
  OAI211_X1 U380 ( .C1(n589), .C2(n163), .A(n164), .B(n165), .ZN(n161) );
  NOR2_X1 U381 ( .A1(A[46]), .A2(B[46]), .ZN(n166) );
  OAI211_X1 U382 ( .C1(A[24]), .C2(B[24]), .A(n326), .B(n325), .ZN(n36) );
  NAND2_X1 U383 ( .A1(A[43]), .A2(B[43]), .ZN(n216) );
  NAND2_X1 U384 ( .A1(A[26]), .A2(B[26]), .ZN(n306) );
  NAND2_X1 U385 ( .A1(B[46]), .A2(A[46]), .ZN(n164) );
  NAND2_X1 U386 ( .A1(B[32]), .A2(A[32]), .ZN(n283) );
  NAND2_X1 U388 ( .A1(B[48]), .A2(A[48]), .ZN(net492609) );
  NOR2_X1 U389 ( .A1(B[40]), .A2(A[40]), .ZN(n77) );
  NAND2_X1 U390 ( .A1(B[21]), .A2(A[21]), .ZN(n401) );
  NAND2_X1 U392 ( .A1(B[25]), .A2(A[25]), .ZN(n369) );
  OR2_X1 U393 ( .A1(B[23]), .A2(A[23]), .ZN(n328) );
  NAND2_X1 U395 ( .A1(A[22]), .A2(B[22]), .ZN(n388) );
  OR2_X1 U396 ( .A1(A[26]), .A2(B[26]), .ZN(n366) );
  NAND2_X1 U397 ( .A1(B[34]), .A2(A[34]), .ZN(n285) );
  NAND2_X1 U398 ( .A1(B[58]), .A2(A[58]), .ZN(net492527) );
  NAND2_X1 U399 ( .A1(B[54]), .A2(A[54]), .ZN(net492568) );
  NAND2_X1 U400 ( .A1(B[40]), .A2(A[40]), .ZN(n222) );
  NAND2_X1 U401 ( .A1(B[50]), .A2(A[50]), .ZN(net492611) );
  OR2_X1 U403 ( .A1(B[24]), .A2(A[24]), .ZN(n372) );
  NAND2_X1 U404 ( .A1(A[18]), .A2(B[18]), .ZN(n428) );
  NAND2_X1 U405 ( .A1(B[23]), .A2(A[23]), .ZN(n399) );
  NAND2_X1 U406 ( .A1(A[19]), .A2(B[19]), .ZN(n414) );
  NAND2_X1 U407 ( .A1(B[62]), .A2(A[62]), .ZN(n120) );
  OR2_X1 U408 ( .A1(B[28]), .A2(A[28]), .ZN(n319) );
  NAND2_X1 U409 ( .A1(A[31]), .A2(B[31]), .ZN(n331) );
  NAND2_X1 U410 ( .A1(B[16]), .A2(A[16]), .ZN(n418) );
  NAND2_X1 U411 ( .A1(A[38]), .A2(B[38]), .ZN(n264) );
  NAND2_X1 U412 ( .A1(A[42]), .A2(B[42]), .ZN(n31) );
  NAND2_X1 U413 ( .A1(A[28]), .A2(B[28]), .ZN(n354) );
  OR2_X1 U414 ( .A1(B[23]), .A2(A[23]), .ZN(n387) );
  NAND2_X1 U415 ( .A1(B[61]), .A2(A[61]), .ZN(n122) );
  OR2_X1 U416 ( .A1(A[40]), .A2(B[40]), .ZN(n79) );
  NAND2_X1 U417 ( .A1(B[63]), .A2(A[63]), .ZN(n119) );
  OR2_X1 U419 ( .A1(A[19]), .A2(B[19]), .ZN(n422) );
  OR2_X1 U420 ( .A1(A[26]), .A2(B[26]), .ZN(n63) );
  OR2_X1 U421 ( .A1(B[61]), .A2(A[61]), .ZN(n133) );
  OR2_X1 U422 ( .A1(A[30]), .A2(B[30]), .ZN(n321) );
  OR2_X1 U423 ( .A1(B[62]), .A2(A[62]), .ZN(n129) );
  OR2_X1 U424 ( .A1(A[31]), .A2(B[31]), .ZN(n322) );
  OR2_X1 U425 ( .A1(B[63]), .A2(A[63]), .ZN(n115) );
  OR2_X1 U426 ( .A1(B[13]), .A2(A[13]), .ZN(n447) );
  OR2_X1 U427 ( .A1(B[14]), .A2(A[14]), .ZN(n445) );
  OR2_X1 U428 ( .A1(B[15]), .A2(A[15]), .ZN(n439) );
  OR2_X1 U429 ( .A1(B[16]), .A2(A[16]), .ZN(n420) );
  INV_X1 U430 ( .A(B[27]), .ZN(n618) );
  OR2_X1 U431 ( .A1(B[6]), .A2(A[6]), .ZN(n106) );
  OR2_X1 U432 ( .A1(B[5]), .A2(A[5]), .ZN(n111) );
  OR2_X1 U433 ( .A1(B[10]), .A2(A[10]), .ZN(n481) );
  OR2_X1 U434 ( .A1(B[9]), .A2(A[9]), .ZN(n93) );
  OR2_X1 U435 ( .A1(B[11]), .A2(A[11]), .ZN(n475) );
  OR2_X1 U436 ( .A1(B[7]), .A2(A[7]), .ZN(n101) );
  OR2_X1 U437 ( .A1(B[8]), .A2(A[8]), .ZN(n97) );
  OR2_X1 U438 ( .A1(B[2]), .A2(A[2]), .ZN(n262) );
  OR2_X1 U439 ( .A1(B[12]), .A2(A[12]), .ZN(n453) );
  OR2_X1 U440 ( .A1(B[1]), .A2(A[1]), .ZN(n350) );
  OR2_X1 U441 ( .A1(B[4]), .A2(A[4]), .ZN(n142) );
  OR2_X1 U442 ( .A1(B[3]), .A2(A[3]), .ZN(n257) );
  OR2_X1 U443 ( .A1(B[0]), .A2(A[0]), .ZN(n494) );
  NAND2_X1 U444 ( .A1(B[14]), .A2(A[14]), .ZN(n443) );
  NAND2_X1 U445 ( .A1(B[1]), .A2(A[1]), .ZN(n349) );
  NAND2_X1 U446 ( .A1(B[8]), .A2(A[8]), .ZN(n98) );
  NAND2_X1 U447 ( .A1(B[12]), .A2(A[12]), .ZN(n450) );
  NAND2_X1 U448 ( .A1(B[6]), .A2(A[6]), .ZN(n103) );
  NAND2_X1 U449 ( .A1(B[13]), .A2(A[13]), .ZN(n449) );
  NAND2_X1 U450 ( .A1(B[9]), .A2(A[9]), .ZN(n94) );
  NAND2_X1 U451 ( .A1(B[2]), .A2(A[2]), .ZN(n259) );
  NAND2_X1 U452 ( .A1(B[0]), .A2(A[0]), .ZN(n425) );
  NAND2_X1 U453 ( .A1(B[4]), .A2(A[4]), .ZN(n141) );
  NAND2_X1 U454 ( .A1(B[5]), .A2(A[5]), .ZN(n110) );
  NAND2_X1 U455 ( .A1(B[10]), .A2(A[10]), .ZN(n478) );
  NAND2_X1 U456 ( .A1(B[3]), .A2(A[3]), .ZN(n258) );
  NAND2_X1 U457 ( .A1(B[7]), .A2(A[7]), .ZN(n102) );
  NAND2_X1 U458 ( .A1(B[15]), .A2(A[15]), .ZN(n441) );
  NAND2_X1 U459 ( .A1(B[11]), .A2(A[11]), .ZN(n479) );
  NOR2_X1 U460 ( .A1(n602), .A2(n68), .ZN(n431) );
  OAI21_X1 U461 ( .B1(n68), .B2(n418), .A(n419), .ZN(n415) );
  INV_X1 U462 ( .A(n68), .ZN(n601) );
  OAI21_X1 U463 ( .B1(n430), .B2(n68), .A(n419), .ZN(n427) );
  NOR2_X1 U464 ( .A1(A[17]), .A2(B[17]), .ZN(n68) );
  NAND2_X1 U465 ( .A1(n245), .A2(n246), .ZN(n192) );
  NAND2_X1 U466 ( .A1(n599), .A2(n246), .ZN(n190) );
  AND2_X1 U467 ( .A1(n246), .A2(n10), .ZN(n84) );
  NAND2_X1 U468 ( .A1(n599), .A2(n246), .ZN(n11) );
  INV_X1 U469 ( .A(net492586), .ZN(n542) );
  NAND2_X1 U470 ( .A1(A[35]), .A2(B[35]), .ZN(n199) );
  OAI22_X1 U471 ( .A1(A[35]), .A2(B[35]), .B1(A[34]), .B2(B[34]), .ZN(n39) );
  XNOR2_X1 U472 ( .A(n375), .B(n32), .ZN(SUM[27]) );
  NAND2_X1 U473 ( .A1(A[47]), .A2(B[47]), .ZN(n158) );
  OAI211_X1 U474 ( .C1(A[47]), .C2(B[47]), .A(n178), .B(n179), .ZN(n176) );
  OR2_X1 U475 ( .A1(A[47]), .A2(B[47]), .ZN(n182) );
  XNOR2_X1 U476 ( .A(n343), .B(n344), .ZN(SUM[30]) );
  INV_X1 U477 ( .A(net492600), .ZN(n571) );
  OR2_X1 U478 ( .A1(A[39]), .A2(B[39]), .ZN(n191) );
  NAND2_X1 U479 ( .A1(B[39]), .A2(A[39]), .ZN(n246) );
  AOI21_X1 U480 ( .B1(n237), .B2(n86), .A(n229), .ZN(n227) );
  NOR2_X1 U481 ( .A1(n594), .A2(n595), .ZN(n228) );
  AOI21_X1 U482 ( .B1(n138), .B2(net492522), .A(n90), .ZN(net492520) );
  AND2_X1 U483 ( .A1(net492533), .A2(net492530), .ZN(n138) );
  AOI21_X1 U484 ( .B1(net537537), .B2(net492604), .A(n585), .ZN(n154) );
  NAND4_X1 U485 ( .A1(n22), .A2(n157), .A3(n158), .A4(n159), .ZN(net537537) );
  NAND2_X1 U486 ( .A1(n160), .A2(n161), .ZN(n159) );
  NAND2_X1 U487 ( .A1(B[36]), .A2(A[36]), .ZN(n249) );
  AOI21_X1 U488 ( .B1(n23), .B2(net492571), .A(n583), .ZN(net492577) );
  NOR2_X1 U489 ( .A1(B[47]), .A2(A[47]), .ZN(n87) );
  OR2_X1 U490 ( .A1(net492559), .A2(n512), .ZN(net538272) );
  NOR2_X1 U491 ( .A1(n580), .A2(n90), .ZN(n144) );
  INV_X1 U492 ( .A(net492533), .ZN(n580) );
  OAI21_X1 U493 ( .B1(n541), .B2(n581), .A(net492526), .ZN(net492546) );
  OAI211_X1 U494 ( .C1(n581), .C2(n51), .A(net492526), .B(net492527), .ZN(
        net492522) );
  NAND2_X1 U495 ( .A1(net492532), .A2(net492526), .ZN(net492553) );
  NAND2_X1 U496 ( .A1(B[57]), .A2(A[57]), .ZN(net492526) );
  OAI211_X1 U497 ( .C1(n282), .C2(n283), .A(n284), .B(n285), .ZN(n281) );
  NAND2_X1 U498 ( .A1(n283), .A2(n284), .ZN(n294) );
  OR2_X1 U499 ( .A1(B[55]), .A2(A[55]), .ZN(net492574) );
  NOR2_X1 U500 ( .A1(n515), .A2(net534634), .ZN(net492578) );
  OAI21_X1 U501 ( .B1(n603), .B2(n323), .A(n562), .ZN(n64) );
  OAI21_X1 U502 ( .B1(n603), .B2(n323), .A(n562), .ZN(n403) );
  AOI21_X1 U503 ( .B1(n249), .B2(n250), .A(n251), .ZN(n248) );
  OAI21_X1 U504 ( .B1(n538), .B2(n575), .A(n120), .ZN(n127) );
  INV_X1 U505 ( .A(n130), .ZN(n538) );
  NOR2_X1 U506 ( .A1(n176), .A2(n177), .ZN(n167) );
  AOI21_X1 U507 ( .B1(n81), .B2(n199), .A(n599), .ZN(n193) );
  AND2_X1 U508 ( .A1(n509), .A2(n81), .ZN(n40) );
  NAND2_X1 U509 ( .A1(n511), .A2(n81), .ZN(n240) );
  INV_X1 U510 ( .A(n115), .ZN(n576) );
  NAND2_X1 U511 ( .A1(n119), .A2(n115), .ZN(n126) );
  XNOR2_X1 U512 ( .A(n130), .B(n131), .ZN(SUM[62]) );
  NAND2_X1 U513 ( .A1(n129), .A2(n120), .ZN(n131) );
  OAI211_X1 U514 ( .C1(n557), .C2(n300), .A(n301), .B(n302), .ZN(n69) );
  NAND2_X1 U515 ( .A1(n179), .A2(n173), .ZN(n297) );
  NAND2_X1 U516 ( .A1(A[30]), .A2(B[30]), .ZN(n332) );
  XNOR2_X1 U517 ( .A(n126), .B(n127), .ZN(SUM[63]) );
  NOR2_X1 U518 ( .A1(B[33]), .A2(A[33]), .ZN(n282) );
  NAND2_X1 U519 ( .A1(B[33]), .A2(A[33]), .ZN(n284) );
  XNOR2_X1 U520 ( .A(n406), .B(n405), .ZN(SUM[23]) );
  NAND2_X1 U521 ( .A1(n388), .A2(n407), .ZN(n406) );
  NAND2_X1 U522 ( .A1(n79), .A2(n518), .ZN(n242) );
  AOI21_X1 U523 ( .B1(n320), .B2(n519), .A(n555), .ZN(n343) );
  NAND2_X1 U524 ( .A1(n357), .A2(n16), .ZN(n355) );
  OAI21_X1 U525 ( .B1(n74), .B2(n589), .A(n165), .ZN(n204) );
  NAND2_X1 U526 ( .A1(B[56]), .A2(A[56]), .ZN(n51) );
  XNOR2_X1 U527 ( .A(n148), .B(n147), .ZN(SUM[51]) );
  XNOR2_X1 U528 ( .A(net538546), .B(net492584), .ZN(SUM[54]) );
  NAND2_X1 U529 ( .A1(B[52]), .A2(A[52]), .ZN(net492566) );
  NAND2_X1 U530 ( .A1(n136), .A2(n123), .ZN(n137) );
  OR2_X1 U531 ( .A1(B[60]), .A2(A[60]), .ZN(n136) );
  OAI21_X1 U532 ( .B1(n594), .B2(n186), .A(n187), .ZN(n184) );
  NAND2_X1 U533 ( .A1(n29), .A2(n186), .ZN(n215) );
  AND2_X1 U534 ( .A1(n186), .A2(n597), .ZN(n86) );
  INV_X1 U535 ( .A(n186), .ZN(n596) );
  NOR2_X1 U536 ( .A1(n87), .A2(n166), .ZN(n160) );
  AND2_X1 U537 ( .A1(net492601), .A2(net492600), .ZN(n47) );
  NAND2_X1 U538 ( .A1(net492608), .A2(net492601), .ZN(n147) );
  NAND4_X1 U539 ( .A1(net492600), .A2(net492601), .A3(n44), .A4(net537537), 
        .ZN(n43) );
  OAI21_X1 U540 ( .B1(n413), .B2(n67), .A(n414), .ZN(n315) );
  NOR2_X1 U541 ( .A1(n329), .A2(n330), .ZN(n300) );
  OAI21_X1 U542 ( .B1(n303), .B2(n13), .A(n89), .ZN(n302) );
  OAI211_X1 U543 ( .C1(n557), .C2(n300), .A(n301), .B(n302), .ZN(n173) );
  OAI21_X1 U544 ( .B1(n50), .B2(n526), .A(net492520), .ZN(net492514) );
  INV_X1 U545 ( .A(net538271), .ZN(n541) );
  OAI21_X1 U546 ( .B1(n526), .B2(n582), .A(n51), .ZN(net538271) );
  XNOR2_X1 U547 ( .A(n263), .B(n84), .ZN(SUM[39]) );
  AOI21_X1 U548 ( .B1(n268), .B2(n252), .A(n598), .ZN(n263) );
  OAI21_X1 U550 ( .B1(n540), .B2(n578), .A(n123), .ZN(n134) );
  OAI21_X1 U551 ( .B1(n540), .B2(n578), .A(n123), .ZN(n21) );
  AOI21_X1 U552 ( .B1(n204), .B2(n169), .A(n591), .ZN(n201) );
  OAI21_X1 U553 ( .B1(n574), .B2(n542), .A(net492567), .ZN(n23) );
  OAI21_X1 U554 ( .B1(n542), .B2(n574), .A(n510), .ZN(net538546) );
  OAI211_X1 U555 ( .C1(n574), .C2(net492566), .A(n510), .B(net492568), .ZN(
        net492563) );
  NAND2_X1 U556 ( .A1(net492573), .A2(net492567), .ZN(net492589) );
  NAND2_X1 U557 ( .A1(A[53]), .A2(B[53]), .ZN(net492567) );
  XNOR2_X1 U558 ( .A(n137), .B(net492514), .ZN(SUM[60]) );
  INV_X1 U559 ( .A(net492514), .ZN(n540) );
  XNOR2_X1 U561 ( .A(n144), .B(n143), .ZN(SUM[59]) );
  NAND2_X1 U562 ( .A1(B[37]), .A2(A[37]), .ZN(n266) );
  NOR2_X1 U564 ( .A1(n248), .A2(n598), .ZN(n245) );
  OR2_X1 U565 ( .A1(A[37]), .A2(B[37]), .ZN(n197) );
  NOR2_X1 U566 ( .A1(A[37]), .A2(B[37]), .ZN(n9) );
  NAND2_X1 U567 ( .A1(A[37]), .A2(B[37]), .ZN(n250) );
  NOR2_X1 U568 ( .A1(B[37]), .A2(A[37]), .ZN(n251) );
  XNOR2_X1 U569 ( .A(n227), .B(n228), .ZN(SUM[43]) );
  NAND2_X1 U571 ( .A1(B[60]), .A2(A[60]), .ZN(n123) );
  XNOR2_X1 U572 ( .A(n134), .B(n135), .ZN(SUM[61]) );
  AND2_X1 U573 ( .A1(n517), .A2(n209), .ZN(n74) );
  AND2_X1 U574 ( .A1(n517), .A2(n209), .ZN(n7) );
  AND2_X1 U575 ( .A1(n152), .A2(n151), .ZN(n71) );
  NAND2_X1 U576 ( .A1(B[49]), .A2(A[49]), .ZN(net492610) );
  OAI211_X1 U577 ( .C1(n540), .C2(n578), .A(n122), .B(n123), .ZN(n117) );
  OAI21_X1 U578 ( .B1(n539), .B2(n577), .A(n122), .ZN(n130) );
  NAND2_X1 U579 ( .A1(n133), .A2(n122), .ZN(n135) );
  AND2_X1 U580 ( .A1(n174), .A2(n172), .ZN(n12) );
  INV_X1 U581 ( .A(n172), .ZN(n588) );
  AND4_X1 U582 ( .A1(n172), .A2(n171), .A3(n568), .A4(n69), .ZN(n88) );
  NOR2_X1 U583 ( .A1(n214), .A2(n587), .ZN(n209) );
  NAND2_X1 U585 ( .A1(n211), .A2(n172), .ZN(n62) );
  NAND2_X1 U586 ( .A1(n172), .A2(n521), .ZN(n217) );
  NAND2_X1 U587 ( .A1(A[44]), .A2(B[44]), .ZN(n163) );
  XNOR2_X1 U588 ( .A(net492577), .B(net492578), .ZN(SUM[55]) );
  NAND2_X1 U590 ( .A1(A[51]), .A2(B[51]), .ZN(net492608) );
  NAND2_X1 U591 ( .A1(n280), .A2(n281), .ZN(n81) );
  NAND2_X1 U592 ( .A1(n280), .A2(n281), .ZN(n198) );
  AOI21_X1 U593 ( .B1(n41), .B2(net492563), .A(net534634), .ZN(net492561) );
  XNOR2_X1 U596 ( .A(net492558), .B(net492555), .ZN(SUM[56]) );
  NAND2_X1 U597 ( .A1(n253), .A2(n249), .ZN(n276) );
  NAND4_X1 U598 ( .A1(n191), .A2(n253), .A3(n197), .A4(n252), .ZN(n175) );
  NAND2_X1 U599 ( .A1(n240), .A2(n253), .ZN(n275) );
  NAND2_X1 U600 ( .A1(n197), .A2(n253), .ZN(n78) );
  INV_X1 U601 ( .A(n253), .ZN(n593) );
  NAND2_X1 U602 ( .A1(n544), .A2(n315), .ZN(n312) );
  XNOR2_X1 U603 ( .A(n408), .B(n409), .ZN(SUM[22]) );
  NAND2_X1 U604 ( .A1(n327), .A2(n408), .ZN(n407) );
  INV_X1 U605 ( .A(n315), .ZN(n562) );
  NAND2_X1 U606 ( .A1(A[17]), .A2(B[17]), .ZN(n419) );
  XNOR2_X1 U607 ( .A(n145), .B(n505), .ZN(SUM[58]) );
  AOI21_X1 U608 ( .B1(net492530), .B2(net492546), .A(n579), .ZN(n143) );
  AND2_X1 U609 ( .A1(B[59]), .A2(A[59]), .ZN(n90) );
  AOI21_X1 U610 ( .B1(n585), .B2(net492625), .A(n572), .ZN(n151) );
  INV_X1 U611 ( .A(net492610), .ZN(n572) );
  XNOR2_X1 U612 ( .A(net538271), .B(net492553), .ZN(SUM[57]) );
  NAND2_X1 U613 ( .A1(net538272), .A2(net492561), .ZN(net492555) );
  AND2_X1 U614 ( .A1(B[55]), .A2(A[55]), .ZN(net534634) );
endmodule


module RCA_NBIT64_8 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_8_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_7_DW01_add_6 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net503772, net503770, net503760, net503756, net503754, net503753,
         net503751, net503748, net503747, net503746, net503732, net503708,
         net503704, net503696, net534635, net536100, net538470, net538671,
         net534627, net503706, net534734, n2, n4, n5, n6, n7, n8, n9, n11, n14,
         n16, n17, n18, n19, n20, n22, n26, n29, n30, n31, n33, n34, n35, n36,
         n37, n38, n41, n42, n44, n45, n48, n49, n50, n51, n52, n53, n55, n57,
         n58, n60, n61, n64, n65, n66, n67, n69, n70, n72, n73, n74, n75, n76,
         n78, n79, n80, n83, n85, n86, n87, n88, n89, n90, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n148, n150, n153, n155, n156, n157, n159, n160, n161,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n188, n189, n190, n191, n193, n194, n195, n196, n197, n199,
         n200, n201, n202, n204, n205, n206, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n244, n245, n246, n249, n250,
         n251, n252, n253, n254, n255, n259, n260, n261, n262, n263, n265,
         n266, n267, n268, n269, n271, n272, n275, n276, n277, n278, n279,
         n280, n282, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n318, n319, n320, n321, n322, n323, n324, n326, n327, n328,
         n329, n331, n332, n335, n338, n339, n340, n341, n343, n344, n345,
         n346, n347, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n364, n365, n367, n368, n371, n372, n373,
         n374, n375, n376, n379, n380, n381, n384, n386, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n409, n410, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n433, n434, n436, n437, n438, n439, n440,
         n441, n443, n445, n446, n447, n448, n449, n452, n453, n454, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n488, n489, n490, n491, n493,
         n494, n495, n496, n497, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602;

  NAND3_X1 U16 ( .A1(n372), .A2(n376), .A3(n5), .ZN(n341) );
  OR2_X2 U61 ( .A1(B[54]), .A2(A[54]), .ZN(net503751) );
  XOR2_X1 U68 ( .A(n410), .B(n510), .Z(SUM[20]) );
  AND2_X2 U105 ( .A1(n51), .A2(n57), .ZN(n58) );
  OR2_X2 U132 ( .A1(B[33]), .A2(A[33]), .ZN(n222) );
  OR2_X2 U388 ( .A1(A[41]), .A2(B[41]), .ZN(n239) );
  NAND3_X1 U509 ( .A1(net503696), .A2(n533), .A3(n157), .ZN(n156) );
  NAND3_X1 U527 ( .A1(n195), .A2(n194), .A3(n196), .ZN(n172) );
  NAND3_X1 U547 ( .A1(n304), .A2(n305), .A3(n306), .ZN(n302) );
  NAND3_X1 U551 ( .A1(n296), .A2(n315), .A3(n316), .ZN(n314) );
  NAND3_X1 U552 ( .A1(n222), .A2(n221), .A3(n213), .ZN(n316) );
  NAND3_X1 U554 ( .A1(n310), .A2(n311), .A3(n312), .ZN(n324) );
  NAND3_X1 U558 ( .A1(n581), .A2(n536), .A3(n538), .ZN(n347) );
  OR2_X2 U134 ( .A1(B[40]), .A2(A[40]), .ZN(n240) );
  OR2_X2 U166 ( .A1(B[46]), .A2(A[46]), .ZN(n212) );
  OR2_X2 U266 ( .A1(B[50]), .A2(A[50]), .ZN(n175) );
  OR2_X2 U371 ( .A1(B[48]), .A2(A[48]), .ZN(n178) );
  OR2_X2 U383 ( .A1(B[32]), .A2(A[32]), .ZN(n221) );
  OR2_X2 U384 ( .A1(B[36]), .A2(A[36]), .ZN(n261) );
  AND2_X1 U2 ( .A1(n493), .A2(n426), .ZN(SUM[0]) );
  OR2_X1 U3 ( .A1(B[58]), .A2(A[58]), .ZN(n160) );
  NOR2_X1 U4 ( .A1(B[61]), .A2(A[61]), .ZN(n521) );
  INV_X1 U5 ( .A(n521), .ZN(n134) );
  INV_X1 U6 ( .A(n522), .ZN(n137) );
  CLKBUF_X1 U7 ( .A(A[51]), .Z(n501) );
  CLKBUF_X1 U8 ( .A(A[30]), .Z(n502) );
  AND2_X1 U9 ( .A1(n554), .A2(net503753), .ZN(n503) );
  OAI211_X1 U10 ( .C1(n266), .C2(n267), .A(n268), .B(n269), .ZN(n504) );
  AOI21_X1 U11 ( .B1(n172), .B2(n178), .A(n556), .ZN(n505) );
  CLKBUF_X1 U12 ( .A(n368), .Z(n506) );
  AOI22_X1 U13 ( .A1(n516), .A2(B[39]), .B1(n571), .B2(n504), .ZN(n507) );
  OAI21_X1 U14 ( .B1(n202), .B2(n75), .A(n199), .ZN(n508) );
  INV_X1 U15 ( .A(n548), .ZN(n509) );
  CLKBUF_X1 U17 ( .A(n70), .Z(n510) );
  NAND3_X1 U18 ( .A1(net503754), .A2(net503751), .A3(n503), .ZN(n50) );
  OAI21_X1 U19 ( .B1(n34), .B2(net536100), .A(net503746), .ZN(n511) );
  OR2_X1 U20 ( .A1(B[53]), .A2(A[53]), .ZN(net503753) );
  OR2_X2 U21 ( .A1(A[25]), .A2(B[25]), .ZN(n375) );
  OR2_X2 U22 ( .A1(A[27]), .A2(B[27]), .ZN(n372) );
  NOR2_X1 U23 ( .A1(A[29]), .A2(B[29]), .ZN(n512) );
  OR2_X1 U24 ( .A1(A[29]), .A2(B[29]), .ZN(n326) );
  NAND3_X1 U25 ( .A1(n195), .A2(n194), .A3(n196), .ZN(n513) );
  AND3_X1 U26 ( .A1(n220), .A2(n212), .A3(n519), .ZN(n514) );
  OR2_X1 U27 ( .A1(A[19]), .A2(B[19]), .ZN(n515) );
  NOR2_X1 U28 ( .A1(B[49]), .A2(A[49]), .ZN(n98) );
  OR2_X1 U29 ( .A1(A[19]), .A2(B[19]), .ZN(n416) );
  CLKBUF_X1 U30 ( .A(A[39]), .Z(n516) );
  OAI21_X1 U31 ( .B1(n232), .B2(n231), .A(n86), .ZN(n517) );
  XNOR2_X1 U32 ( .A(n244), .B(n518), .ZN(SUM[43]) );
  NAND2_X1 U33 ( .A1(n86), .A2(n234), .ZN(n518) );
  AND2_X1 U34 ( .A1(n219), .A2(n218), .ZN(n519) );
  AND3_X1 U35 ( .A1(n220), .A2(n212), .A3(n519), .ZN(n96) );
  OR2_X1 U36 ( .A1(B[44]), .A2(A[44]), .ZN(n218) );
  OR2_X1 U37 ( .A1(B[42]), .A2(A[42]), .ZN(n241) );
  NAND4_X2 U38 ( .A1(n305), .A2(n307), .A3(n322), .A4(n308), .ZN(n213) );
  CLKBUF_X1 U39 ( .A(net536100), .Z(n520) );
  AND2_X1 U40 ( .A1(n171), .A2(n170), .ZN(net536100) );
  AND2_X2 U41 ( .A1(n156), .A2(n155), .ZN(n522) );
  NOR2_X1 U42 ( .A1(A[57]), .A2(B[57]), .ZN(net534734) );
  XOR2_X1 U43 ( .A(n90), .B(n523), .Z(SUM[35]) );
  NAND2_X1 U44 ( .A1(n217), .A2(n297), .ZN(n523) );
  XOR2_X1 U45 ( .A(n524), .B(n242), .Z(SUM[40]) );
  AND2_X1 U46 ( .A1(n240), .A2(n253), .ZN(n524) );
  NOR2_X1 U47 ( .A1(n79), .A2(n343), .ZN(n70) );
  NOR2_X1 U48 ( .A1(n585), .A2(n351), .ZN(n79) );
  NOR2_X1 U49 ( .A1(n204), .A2(n575), .ZN(n286) );
  INV_X1 U50 ( .A(A[31]), .ZN(n579) );
  INV_X1 U51 ( .A(n350), .ZN(n536) );
  NAND2_X1 U52 ( .A1(n536), .A2(n343), .ZN(n340) );
  INV_X1 U53 ( .A(n58), .ZN(n533) );
  OAI21_X1 U54 ( .B1(n598), .B2(n461), .A(n458), .ZN(n109) );
  AOI21_X1 U55 ( .B1(n457), .B2(n458), .A(n459), .ZN(n454) );
  NAND2_X1 U56 ( .A1(n593), .A2(n460), .ZN(n457) );
  INV_X1 U57 ( .A(n461), .ZN(n593) );
  NAND2_X1 U58 ( .A1(n473), .A2(n456), .ZN(n471) );
  NAND2_X1 U59 ( .A1(n590), .A2(n109), .ZN(n473) );
  INV_X1 U60 ( .A(n459), .ZN(n590) );
  INV_X1 U62 ( .A(n460), .ZN(n598) );
  INV_X1 U63 ( .A(n344), .ZN(n585) );
  INV_X1 U64 ( .A(n341), .ZN(n538) );
  INV_X1 U65 ( .A(n351), .ZN(n581) );
  INV_X1 U66 ( .A(n456), .ZN(n589) );
  INV_X1 U67 ( .A(n126), .ZN(SUM[64]) );
  NAND2_X1 U69 ( .A1(n181), .A2(n178), .ZN(n193) );
  AND2_X1 U70 ( .A1(n259), .A2(n66), .ZN(n75) );
  NOR2_X1 U71 ( .A1(n94), .A2(n99), .ZN(n66) );
  NAND2_X1 U72 ( .A1(n401), .A2(n400), .ZN(n410) );
  NOR2_X1 U73 ( .A1(n565), .A2(n566), .ZN(n255) );
  AOI21_X1 U74 ( .B1(n242), .B2(n240), .A(n238), .ZN(n254) );
  INV_X1 U75 ( .A(n239), .ZN(n566) );
  AND3_X1 U76 ( .A1(n396), .A2(n397), .A3(n398), .ZN(n17) );
  NAND2_X1 U77 ( .A1(n399), .A2(n400), .ZN(n397) );
  INV_X1 U78 ( .A(n31), .ZN(n539) );
  NAND2_X1 U79 ( .A1(n597), .A2(n579), .ZN(n331) );
  NAND2_X1 U80 ( .A1(n221), .A2(n294), .ZN(n321) );
  NOR2_X1 U81 ( .A1(n99), .A2(n572), .ZN(n88) );
  NOR2_X1 U82 ( .A1(n555), .A2(n34), .ZN(net503772) );
  INV_X1 U83 ( .A(net503746), .ZN(n555) );
  NAND2_X1 U84 ( .A1(n379), .A2(n578), .ZN(n391) );
  NAND2_X1 U85 ( .A1(n267), .A2(n261), .ZN(n285) );
  NAND2_X1 U86 ( .A1(n296), .A2(n222), .ZN(n318) );
  NAND2_X1 U87 ( .A1(n367), .A2(n327), .ZN(n89) );
  NAND2_X1 U88 ( .A1(n398), .A2(n395), .ZN(n406) );
  INV_X1 U89 ( .A(net503748), .ZN(n552) );
  NOR2_X1 U90 ( .A1(n558), .A2(n98), .ZN(n191) );
  INV_X1 U91 ( .A(n182), .ZN(n558) );
  NAND2_X1 U92 ( .A1(n396), .A2(n399), .ZN(n409) );
  NAND2_X1 U93 ( .A1(n263), .A2(n268), .ZN(n282) );
  INV_X1 U94 ( .A(n181), .ZN(n556) );
  NAND2_X1 U95 ( .A1(net503751), .A2(net503748), .ZN(n169) );
  NAND2_X1 U96 ( .A1(n218), .A2(n208), .ZN(n230) );
  NAND2_X1 U97 ( .A1(n175), .A2(n183), .ZN(n188) );
  NAND2_X1 U98 ( .A1(n212), .A2(n210), .ZN(n228) );
  AND2_X1 U99 ( .A1(n375), .A2(n379), .ZN(n5) );
  NAND2_X1 U100 ( .A1(n323), .A2(n324), .ZN(n322) );
  NOR2_X1 U101 ( .A1(n328), .A2(n26), .ZN(n323) );
  XNOR2_X1 U102 ( .A(n380), .B(n381), .ZN(SUM[27]) );
  NOR2_X1 U103 ( .A1(n545), .A2(n544), .ZN(n381) );
  AOI21_X1 U104 ( .B1(n384), .B2(n376), .A(n541), .ZN(n380) );
  INV_X1 U106 ( .A(n373), .ZN(n545) );
  OAI21_X1 U107 ( .B1(n74), .B2(n543), .A(n542), .ZN(n384) );
  INV_X1 U108 ( .A(n375), .ZN(n543) );
  XNOR2_X1 U109 ( .A(n384), .B(n386), .ZN(SUM[26]) );
  NAND2_X1 U110 ( .A1(n376), .A2(n374), .ZN(n386) );
  OAI21_X1 U111 ( .B1(n413), .B2(n412), .A(n414), .ZN(n343) );
  NOR2_X1 U112 ( .A1(n417), .A2(n418), .ZN(n412) );
  NAND2_X1 U113 ( .A1(n416), .A2(n415), .ZN(n413) );
  NOR2_X1 U114 ( .A1(n582), .A2(n422), .ZN(n417) );
  AND2_X1 U115 ( .A1(n219), .A2(n209), .ZN(n8) );
  NAND2_X1 U116 ( .A1(n239), .A2(n241), .ZN(n245) );
  AOI21_X1 U117 ( .B1(n291), .B2(n315), .A(n292), .ZN(n204) );
  AND2_X1 U118 ( .A1(n295), .A2(n296), .ZN(n291) );
  NAND2_X1 U119 ( .A1(n293), .A2(n69), .ZN(n292) );
  INV_X1 U120 ( .A(net503708), .ZN(n547) );
  NOR2_X1 U121 ( .A1(n569), .A2(n101), .ZN(n225) );
  INV_X1 U122 ( .A(n220), .ZN(n569) );
  NAND2_X1 U123 ( .A1(n326), .A2(n576), .ZN(n310) );
  INV_X1 U124 ( .A(n327), .ZN(n576) );
  XNOR2_X1 U125 ( .A(n355), .B(n356), .ZN(SUM[30]) );
  NAND2_X1 U126 ( .A1(n335), .A2(n312), .ZN(n356) );
  NAND2_X1 U127 ( .A1(n223), .A2(n222), .ZN(n301) );
  AOI21_X1 U128 ( .B1(n302), .B2(n221), .A(n303), .ZN(n300) );
  NAND2_X1 U129 ( .A1(n294), .A2(n296), .ZN(n303) );
  XNOR2_X1 U130 ( .A(n141), .B(n142), .ZN(SUM[63]) );
  NAND2_X1 U131 ( .A1(n130), .A2(n129), .ZN(n141) );
  NAND2_X1 U133 ( .A1(n135), .A2(n144), .ZN(n143) );
  XNOR2_X1 U135 ( .A(n358), .B(n365), .ZN(SUM[29]) );
  NAND2_X1 U136 ( .A1(n326), .A2(n311), .ZN(n365) );
  OAI21_X1 U137 ( .B1(n529), .B2(n577), .A(n327), .ZN(n358) );
  NOR2_X1 U138 ( .A1(n299), .A2(n574), .ZN(n90) );
  INV_X1 U139 ( .A(n295), .ZN(n574) );
  OAI21_X1 U140 ( .B1(n341), .B2(n530), .A(n338), .ZN(n368) );
  OAI21_X1 U141 ( .B1(n540), .B2(n371), .A(n372), .ZN(n338) );
  NAND2_X1 U142 ( .A1(n234), .A2(n235), .ZN(n232) );
  NAND2_X1 U143 ( .A1(n238), .A2(n239), .ZN(n236) );
  INV_X1 U144 ( .A(n33), .ZN(n549) );
  OAI211_X1 U145 ( .C1(n98), .C2(n181), .A(n182), .B(n183), .ZN(n180) );
  XNOR2_X1 U146 ( .A(n388), .B(n389), .ZN(SUM[25]) );
  NAND2_X1 U147 ( .A1(n375), .A2(n542), .ZN(n389) );
  NAND2_X1 U148 ( .A1(n390), .A2(n578), .ZN(n388) );
  XNOR2_X1 U149 ( .A(n403), .B(n402), .ZN(SUM[23]) );
  INV_X1 U150 ( .A(n367), .ZN(n577) );
  XNOR2_X1 U151 ( .A(n313), .B(n314), .ZN(SUM[34]) );
  NAND2_X1 U152 ( .A1(n223), .A2(n295), .ZN(n313) );
  AND2_X1 U153 ( .A1(n525), .A2(n262), .ZN(n284) );
  AOI21_X1 U154 ( .B1(n261), .B2(n260), .A(n93), .ZN(n61) );
  OAI21_X1 U155 ( .B1(n540), .B2(n371), .A(n372), .ZN(n31) );
  OR2_X1 U156 ( .A1(n197), .A2(n563), .ZN(n87) );
  AOI21_X1 U157 ( .B1(n200), .B2(n201), .A(n202), .ZN(n197) );
  OAI21_X1 U158 ( .B1(n562), .B2(n11), .A(n240), .ZN(n7) );
  AOI21_X1 U159 ( .B1(n565), .B2(n241), .A(n564), .ZN(n246) );
  INV_X1 U160 ( .A(net503751), .ZN(n553) );
  NOR2_X1 U161 ( .A1(n289), .A2(n290), .ZN(n288) );
  NAND2_X1 U162 ( .A1(n69), .A2(n222), .ZN(n290) );
  NAND2_X1 U163 ( .A1(n217), .A2(n221), .ZN(n289) );
  OAI211_X1 U164 ( .C1(n551), .C2(net503746), .A(net503747), .B(net503748), 
        .ZN(n53) );
  NOR2_X1 U165 ( .A1(n99), .A2(n94), .ZN(n200) );
  NAND2_X1 U167 ( .A1(n309), .A2(n324), .ZN(n304) );
  AND2_X1 U168 ( .A1(n307), .A2(n308), .ZN(n306) );
  NOR2_X1 U169 ( .A1(n328), .A2(n26), .ZN(n309) );
  INV_X1 U170 ( .A(n237), .ZN(n565) );
  NAND2_X1 U171 ( .A1(n357), .A2(n311), .ZN(n355) );
  OAI21_X1 U172 ( .B1(n529), .B2(n577), .A(n327), .ZN(n65) );
  NAND2_X1 U173 ( .A1(n373), .A2(n374), .ZN(n371) );
  NAND2_X1 U174 ( .A1(n393), .A2(n16), .ZN(n350) );
  AND3_X1 U175 ( .A1(n398), .A2(n396), .A3(n401), .ZN(n16) );
  OAI21_X1 U176 ( .B1(n11), .B2(n562), .A(n240), .ZN(n252) );
  AOI21_X1 U177 ( .B1(net503732), .B2(n548), .A(n33), .ZN(n41) );
  NAND2_X1 U178 ( .A1(n560), .A2(n222), .ZN(n315) );
  INV_X1 U179 ( .A(n294), .ZN(n560) );
  NOR2_X1 U180 ( .A1(n98), .A2(n557), .ZN(n174) );
  INV_X1 U181 ( .A(n178), .ZN(n557) );
  INV_X1 U182 ( .A(n36), .ZN(n578) );
  NAND2_X1 U183 ( .A1(n419), .A2(n420), .ZN(n418) );
  AOI21_X1 U184 ( .B1(n179), .B2(n180), .A(n97), .ZN(n170) );
  AND3_X1 U185 ( .A1(n176), .A2(n174), .A3(n175), .ZN(n173) );
  INV_X1 U186 ( .A(n37), .ZN(n542) );
  INV_X1 U187 ( .A(n235), .ZN(n564) );
  INV_X1 U188 ( .A(n297), .ZN(n575) );
  AOI21_X1 U189 ( .B1(n249), .B2(n239), .A(n565), .ZN(n250) );
  NAND2_X1 U190 ( .A1(n7), .A2(n253), .ZN(n249) );
  NAND2_X1 U191 ( .A1(n76), .A2(n217), .ZN(n216) );
  INV_X1 U192 ( .A(n374), .ZN(n541) );
  INV_X1 U193 ( .A(n208), .ZN(n570) );
  INV_X1 U194 ( .A(n262), .ZN(n561) );
  AND2_X1 U195 ( .A1(n176), .A2(n175), .ZN(n179) );
  INV_X1 U196 ( .A(n396), .ZN(n537) );
  INV_X1 U197 ( .A(n372), .ZN(n544) );
  INV_X1 U198 ( .A(n528), .ZN(n139) );
  INV_X1 U199 ( .A(n268), .ZN(n573) );
  AND2_X1 U200 ( .A1(n215), .A2(n18), .ZN(n6) );
  NOR2_X1 U201 ( .A1(n202), .A2(n216), .ZN(n215) );
  AND3_X1 U202 ( .A1(n223), .A2(n222), .A3(n221), .ZN(n214) );
  AND2_X1 U203 ( .A1(n29), .A2(n212), .ZN(n205) );
  INV_X1 U204 ( .A(n183), .ZN(n559) );
  INV_X1 U205 ( .A(n210), .ZN(n568) );
  XNOR2_X1 U206 ( .A(n427), .B(n428), .ZN(SUM[19]) );
  NAND2_X1 U207 ( .A1(n419), .A2(n429), .ZN(n428) );
  NAND2_X1 U208 ( .A1(n515), .A2(n414), .ZN(n427) );
  NAND2_X1 U209 ( .A1(n415), .A2(n430), .ZN(n429) );
  XNOR2_X1 U210 ( .A(n462), .B(n463), .ZN(SUM[15]) );
  NAND2_X1 U211 ( .A1(n464), .A2(n447), .ZN(n463) );
  NAND2_X1 U212 ( .A1(n443), .A2(n449), .ZN(n462) );
  NAND2_X1 U213 ( .A1(n448), .A2(n465), .ZN(n464) );
  XNOR2_X1 U214 ( .A(n431), .B(n430), .ZN(SUM[18]) );
  NAND2_X1 U215 ( .A1(n415), .A2(n419), .ZN(n431) );
  XNOR2_X1 U216 ( .A(n466), .B(n465), .ZN(SUM[14]) );
  NAND2_X1 U217 ( .A1(n448), .A2(n447), .ZN(n466) );
  XNOR2_X1 U218 ( .A(n434), .B(n433), .ZN(SUM[17]) );
  NAND2_X1 U219 ( .A1(n424), .A2(n420), .ZN(n434) );
  XNOR2_X1 U220 ( .A(n469), .B(n468), .ZN(SUM[13]) );
  NAND2_X1 U221 ( .A1(n453), .A2(n446), .ZN(n469) );
  XNOR2_X1 U222 ( .A(n436), .B(n344), .ZN(SUM[16]) );
  NAND2_X1 U223 ( .A1(n423), .A2(n422), .ZN(n436) );
  XNOR2_X1 U224 ( .A(n112), .B(n113), .ZN(SUM[7]) );
  NAND2_X1 U225 ( .A1(n116), .A2(n117), .ZN(n112) );
  NAND2_X1 U226 ( .A1(n114), .A2(n115), .ZN(n113) );
  NAND2_X1 U227 ( .A1(n118), .A2(n119), .ZN(n117) );
  XNOR2_X1 U228 ( .A(n271), .B(n272), .ZN(SUM[3]) );
  OAI21_X1 U229 ( .B1(n601), .B2(n599), .A(n275), .ZN(n272) );
  NAND2_X1 U230 ( .A1(n277), .A2(n278), .ZN(n271) );
  INV_X1 U231 ( .A(n276), .ZN(n601) );
  XNOR2_X1 U232 ( .A(n425), .B(n602), .ZN(SUM[1]) );
  NAND2_X1 U233 ( .A1(n362), .A2(n361), .ZN(n425) );
  XNOR2_X1 U234 ( .A(n472), .B(n471), .ZN(SUM[12]) );
  NAND2_X1 U235 ( .A1(n452), .A2(n445), .ZN(n472) );
  XNOR2_X1 U236 ( .A(n108), .B(n109), .ZN(SUM[8]) );
  NAND2_X1 U237 ( .A1(n110), .A2(n111), .ZN(n108) );
  XNOR2_X1 U238 ( .A(n359), .B(n276), .ZN(SUM[2]) );
  NAND2_X1 U239 ( .A1(n364), .A2(n275), .ZN(n359) );
  XNOR2_X1 U240 ( .A(n161), .B(n125), .ZN(SUM[5]) );
  NAND2_X1 U241 ( .A1(n124), .A2(n123), .ZN(n161) );
  XNOR2_X1 U242 ( .A(n485), .B(n484), .ZN(SUM[10]) );
  NAND2_X1 U243 ( .A1(n480), .A2(n478), .ZN(n485) );
  XNOR2_X1 U244 ( .A(n481), .B(n482), .ZN(SUM[11]) );
  NAND2_X1 U245 ( .A1(n478), .A2(n483), .ZN(n482) );
  NAND2_X1 U246 ( .A1(n477), .A2(n476), .ZN(n481) );
  NAND2_X1 U247 ( .A1(n480), .A2(n484), .ZN(n483) );
  XNOR2_X1 U248 ( .A(n120), .B(n118), .ZN(SUM[6]) );
  NAND2_X1 U249 ( .A1(n119), .A2(n116), .ZN(n120) );
  XNOR2_X1 U250 ( .A(n104), .B(n105), .ZN(SUM[9]) );
  NAND2_X1 U251 ( .A1(n106), .A2(n107), .ZN(n104) );
  XNOR2_X1 U252 ( .A(n190), .B(n460), .ZN(SUM[4]) );
  NAND2_X1 U253 ( .A1(n164), .A2(n163), .ZN(n190) );
  OAI21_X1 U254 ( .B1(n494), .B2(n495), .A(n278), .ZN(n460) );
  NAND2_X1 U255 ( .A1(n364), .A2(n277), .ZN(n495) );
  NOR2_X1 U256 ( .A1(n496), .A2(n497), .ZN(n494) );
  NAND2_X1 U257 ( .A1(n275), .A2(n361), .ZN(n497) );
  OAI21_X1 U258 ( .B1(n437), .B2(n438), .A(n439), .ZN(n344) );
  NOR2_X1 U259 ( .A1(n454), .A2(n589), .ZN(n437) );
  NAND4_X1 U260 ( .A1(n452), .A2(n453), .A3(n448), .A4(n449), .ZN(n438) );
  AOI21_X1 U261 ( .B1(n440), .B2(n441), .A(n586), .ZN(n439) );
  OAI21_X1 U262 ( .B1(n592), .B2(n591), .A(n107), .ZN(n484) );
  INV_X1 U263 ( .A(n105), .ZN(n592) );
  INV_X1 U264 ( .A(n106), .ZN(n591) );
  OAI21_X1 U265 ( .B1(n588), .B2(n587), .A(n446), .ZN(n465) );
  INV_X1 U267 ( .A(n468), .ZN(n588) );
  OAI21_X1 U268 ( .B1(n583), .B2(n582), .A(n420), .ZN(n430) );
  INV_X1 U269 ( .A(n433), .ZN(n583) );
  OAI21_X1 U270 ( .B1(n585), .B2(n584), .A(n422), .ZN(n433) );
  INV_X1 U271 ( .A(n423), .ZN(n584) );
  OAI21_X1 U272 ( .B1(n596), .B2(n598), .A(n163), .ZN(n125) );
  INV_X1 U273 ( .A(n164), .ZN(n596) );
  NAND2_X1 U274 ( .A1(n139), .A2(n140), .ZN(n138) );
  OAI21_X1 U275 ( .B1(n595), .B2(n594), .A(n123), .ZN(n118) );
  INV_X1 U276 ( .A(n125), .ZN(n595) );
  INV_X1 U277 ( .A(n124), .ZN(n594) );
  OAI21_X1 U278 ( .B1(n474), .B2(n475), .A(n476), .ZN(n456) );
  NAND2_X1 U279 ( .A1(n477), .A2(n478), .ZN(n475) );
  NOR2_X1 U280 ( .A1(n19), .A2(n479), .ZN(n474) );
  AND2_X1 U281 ( .A1(n107), .A2(n111), .ZN(n19) );
  OAI21_X1 U282 ( .B1(n489), .B2(n490), .A(n114), .ZN(n458) );
  NAND2_X1 U283 ( .A1(n115), .A2(n116), .ZN(n490) );
  NOR2_X1 U284 ( .A1(n20), .A2(n491), .ZN(n489) );
  AND2_X1 U285 ( .A1(n123), .A2(n163), .ZN(n20) );
  NAND4_X1 U286 ( .A1(n423), .A2(n424), .A3(n415), .A4(n515), .ZN(n351) );
  NAND4_X1 U287 ( .A1(n164), .A2(n124), .A3(n119), .A4(n114), .ZN(n461) );
  NAND4_X1 U288 ( .A1(n106), .A2(n110), .A3(n480), .A4(n476), .ZN(n459) );
  OAI211_X1 U289 ( .C1(n587), .C2(n445), .A(n446), .B(n447), .ZN(n441) );
  NAND4_X1 U290 ( .A1(n335), .A2(n344), .A3(n345), .A4(n346), .ZN(n305) );
  NOR2_X1 U291 ( .A1(n512), .A2(n577), .ZN(n345) );
  NOR2_X1 U292 ( .A1(n347), .A2(n328), .ZN(n346) );
  OAI21_X1 U293 ( .B1(n127), .B2(n128), .A(n129), .ZN(n126) );
  NOR2_X1 U294 ( .A1(n132), .A2(n133), .ZN(n127) );
  NOR2_X1 U295 ( .A1(n600), .A2(n426), .ZN(n496) );
  INV_X1 U296 ( .A(n362), .ZN(n600) );
  NAND2_X1 U297 ( .A1(n360), .A2(n361), .ZN(n276) );
  NAND2_X1 U298 ( .A1(n362), .A2(n602), .ZN(n360) );
  NAND2_X1 U299 ( .A1(n470), .A2(n445), .ZN(n468) );
  NAND2_X1 U300 ( .A1(n471), .A2(n452), .ZN(n470) );
  NAND2_X1 U301 ( .A1(n488), .A2(n111), .ZN(n105) );
  NAND2_X1 U302 ( .A1(n109), .A2(n110), .ZN(n488) );
  INV_X1 U303 ( .A(n426), .ZN(n602) );
  INV_X1 U304 ( .A(n424), .ZN(n582) );
  INV_X1 U305 ( .A(n453), .ZN(n587) );
  NAND2_X1 U306 ( .A1(n124), .A2(n119), .ZN(n491) );
  NAND2_X1 U307 ( .A1(n480), .A2(n106), .ZN(n479) );
  AND2_X1 U308 ( .A1(n449), .A2(n448), .ZN(n440) );
  INV_X1 U309 ( .A(n364), .ZN(n599) );
  INV_X1 U310 ( .A(n443), .ZN(n586) );
  NOR2_X1 U311 ( .A1(A[31]), .A2(B[31]), .ZN(n328) );
  NOR2_X1 U312 ( .A1(n72), .A2(n97), .ZN(n185) );
  NOR2_X1 U313 ( .A1(B[56]), .A2(A[56]), .ZN(net534627) );
  NOR2_X1 U314 ( .A1(B[30]), .A2(A[30]), .ZN(n26) );
  OAI211_X1 U315 ( .C1(n266), .C2(n267), .A(n268), .B(n269), .ZN(n265) );
  NOR3_X1 U316 ( .A1(n78), .A2(n577), .A3(n512), .ZN(n332) );
  NOR2_X1 U317 ( .A1(A[30]), .A2(B[30]), .ZN(n78) );
  NAND2_X1 U318 ( .A1(B[28]), .A2(A[28]), .ZN(n327) );
  OAI21_X1 U319 ( .B1(n70), .B2(n2), .A(n400), .ZN(n42) );
  NOR2_X1 U320 ( .A1(A[20]), .A2(B[20]), .ZN(n2) );
  NAND2_X1 U321 ( .A1(B[32]), .A2(A[32]), .ZN(n294) );
  NAND2_X1 U322 ( .A1(B[26]), .A2(A[26]), .ZN(n374) );
  NAND2_X1 U323 ( .A1(A[20]), .A2(B[20]), .ZN(n400) );
  OR2_X1 U324 ( .A1(B[18]), .A2(A[18]), .ZN(n415) );
  NAND2_X1 U325 ( .A1(B[31]), .A2(A[31]), .ZN(n308) );
  NAND2_X1 U326 ( .A1(A[30]), .A2(B[30]), .ZN(n312) );
  NAND2_X1 U327 ( .A1(B[21]), .A2(A[21]), .ZN(n399) );
  NAND3_X1 U328 ( .A1(n241), .A2(n233), .A3(n73), .ZN(n202) );
  OR2_X1 U329 ( .A1(A[43]), .A2(B[43]), .ZN(n233) );
  AND2_X1 U330 ( .A1(n239), .A2(n240), .ZN(n73) );
  NAND2_X1 U331 ( .A1(B[33]), .A2(A[33]), .ZN(n296) );
  NAND2_X1 U332 ( .A1(B[38]), .A2(A[38]), .ZN(n268) );
  NAND2_X1 U333 ( .A1(B[50]), .A2(A[50]), .ZN(n183) );
  NAND2_X1 U334 ( .A1(A[34]), .A2(B[34]), .ZN(n295) );
  NOR2_X1 U335 ( .A1(A[42]), .A2(B[42]), .ZN(n83) );
  NAND2_X1 U336 ( .A1(A[49]), .A2(B[49]), .ZN(n182) );
  NAND2_X1 U337 ( .A1(B[48]), .A2(A[48]), .ZN(n181) );
  NAND2_X1 U338 ( .A1(A[52]), .A2(B[52]), .ZN(net503746) );
  NAND2_X1 U339 ( .A1(A[29]), .A2(B[29]), .ZN(n311) );
  NAND2_X1 U340 ( .A1(B[40]), .A2(A[40]), .ZN(n253) );
  NAND2_X1 U341 ( .A1(B[46]), .A2(A[46]), .ZN(n210) );
  NAND2_X1 U342 ( .A1(B[44]), .A2(A[44]), .ZN(n208) );
  OR2_X1 U343 ( .A1(A[21]), .A2(B[21]), .ZN(n396) );
  OR2_X1 U344 ( .A1(B[30]), .A2(n502), .ZN(n335) );
  NAND2_X1 U345 ( .A1(n507), .A2(n259), .ZN(n242) );
  NAND2_X1 U346 ( .A1(A[27]), .A2(B[27]), .ZN(n373) );
  AND2_X1 U347 ( .A1(B[24]), .A2(A[24]), .ZN(n36) );
  NAND2_X1 U348 ( .A1(B[22]), .A2(A[22]), .ZN(n395) );
  OR2_X1 U349 ( .A1(B[22]), .A2(A[22]), .ZN(n398) );
  NAND2_X1 U350 ( .A1(B[36]), .A2(A[36]), .ZN(n267) );
  OR2_X1 U351 ( .A1(B[24]), .A2(A[24]), .ZN(n379) );
  INV_X1 U352 ( .A(n34), .ZN(n554) );
  OR2_X1 U353 ( .A1(A[26]), .A2(B[26]), .ZN(n376) );
  OR2_X1 U354 ( .A1(A[34]), .A2(B[34]), .ZN(n223) );
  NAND2_X1 U355 ( .A1(B[62]), .A2(A[62]), .ZN(n131) );
  NAND2_X1 U356 ( .A1(A[23]), .A2(B[23]), .ZN(n394) );
  NAND2_X1 U357 ( .A1(B[41]), .A2(A[41]), .ZN(n237) );
  AND2_X1 U358 ( .A1(B[40]), .A2(A[40]), .ZN(n238) );
  AND2_X1 U359 ( .A1(A[25]), .A2(B[25]), .ZN(n37) );
  OR2_X1 U360 ( .A1(B[23]), .A2(A[23]), .ZN(n393) );
  OR2_X1 U361 ( .A1(A[45]), .A2(B[45]), .ZN(n219) );
  OR2_X1 U362 ( .A1(B[62]), .A2(A[62]), .ZN(n135) );
  OR2_X1 U363 ( .A1(B[38]), .A2(A[38]), .ZN(n263) );
  OR2_X1 U364 ( .A1(B[63]), .A2(A[63]), .ZN(n129) );
  OR2_X1 U365 ( .A1(A[34]), .A2(B[34]), .ZN(n69) );
  INV_X1 U366 ( .A(n45), .ZN(n540) );
  OAI221_X1 U367 ( .B1(B[26]), .B2(A[26]), .C1(n37), .C2(n36), .A(n375), .ZN(
        n45) );
  OR2_X1 U368 ( .A1(A[35]), .A2(B[35]), .ZN(n217) );
  OR2_X1 U369 ( .A1(B[28]), .A2(A[28]), .ZN(n367) );
  AND2_X1 U370 ( .A1(A[47]), .A2(B[47]), .ZN(n101) );
  INV_X1 U372 ( .A(n38), .ZN(n571) );
  AND2_X1 U373 ( .A1(B[36]), .A2(A[36]), .ZN(n93) );
  OR2_X1 U374 ( .A1(A[47]), .A2(B[47]), .ZN(n29) );
  OR2_X1 U375 ( .A1(A[43]), .A2(B[43]), .ZN(n86) );
  OR2_X1 U376 ( .A1(A[20]), .A2(B[20]), .ZN(n401) );
  XNOR2_X1 U377 ( .A(n352), .B(n353), .ZN(SUM[31]) );
  OAI21_X1 U378 ( .B1(A[31]), .B2(B[31]), .A(n308), .ZN(n353) );
  NAND2_X1 U379 ( .A1(n354), .A2(n312), .ZN(n352) );
  NAND2_X1 U380 ( .A1(n355), .A2(n335), .ZN(n354) );
  OR2_X1 U381 ( .A1(B[47]), .A2(A[47]), .ZN(n220) );
  NAND2_X1 U382 ( .A1(A[37]), .A2(B[37]), .ZN(n525) );
  OR2_X1 U385 ( .A1(B[14]), .A2(A[14]), .ZN(n448) );
  OR2_X1 U386 ( .A1(B[17]), .A2(A[17]), .ZN(n424) );
  OR2_X1 U387 ( .A1(B[13]), .A2(A[13]), .ZN(n453) );
  OR2_X1 U389 ( .A1(B[16]), .A2(A[16]), .ZN(n423) );
  OR2_X1 U390 ( .A1(B[15]), .A2(A[15]), .ZN(n449) );
  INV_X1 U391 ( .A(B[31]), .ZN(n597) );
  OR2_X1 U392 ( .A1(B[6]), .A2(A[6]), .ZN(n119) );
  OR2_X1 U393 ( .A1(B[9]), .A2(A[9]), .ZN(n106) );
  OR2_X1 U394 ( .A1(B[10]), .A2(A[10]), .ZN(n480) );
  OR2_X1 U395 ( .A1(B[5]), .A2(A[5]), .ZN(n124) );
  OR2_X1 U396 ( .A1(B[11]), .A2(A[11]), .ZN(n476) );
  OR2_X1 U397 ( .A1(B[7]), .A2(A[7]), .ZN(n114) );
  OR2_X1 U398 ( .A1(B[8]), .A2(A[8]), .ZN(n110) );
  OR2_X1 U399 ( .A1(B[12]), .A2(A[12]), .ZN(n452) );
  OR2_X1 U400 ( .A1(B[1]), .A2(A[1]), .ZN(n362) );
  OR2_X1 U401 ( .A1(B[2]), .A2(A[2]), .ZN(n364) );
  OR2_X1 U402 ( .A1(B[4]), .A2(A[4]), .ZN(n164) );
  OR2_X1 U403 ( .A1(B[3]), .A2(A[3]), .ZN(n277) );
  OR2_X1 U404 ( .A1(B[0]), .A2(A[0]), .ZN(n493) );
  NAND2_X1 U405 ( .A1(B[1]), .A2(A[1]), .ZN(n361) );
  NAND2_X1 U406 ( .A1(B[17]), .A2(A[17]), .ZN(n420) );
  NAND2_X1 U407 ( .A1(B[12]), .A2(A[12]), .ZN(n445) );
  NAND2_X1 U408 ( .A1(B[14]), .A2(A[14]), .ZN(n447) );
  NAND2_X1 U409 ( .A1(B[16]), .A2(A[16]), .ZN(n422) );
  NAND2_X1 U410 ( .A1(B[13]), .A2(A[13]), .ZN(n446) );
  NAND2_X1 U411 ( .A1(B[6]), .A2(A[6]), .ZN(n116) );
  NAND2_X1 U412 ( .A1(B[10]), .A2(A[10]), .ZN(n478) );
  NAND2_X1 U413 ( .A1(B[2]), .A2(A[2]), .ZN(n275) );
  NAND2_X1 U414 ( .A1(B[8]), .A2(A[8]), .ZN(n111) );
  NAND2_X1 U415 ( .A1(B[0]), .A2(A[0]), .ZN(n426) );
  NAND2_X1 U416 ( .A1(B[4]), .A2(A[4]), .ZN(n163) );
  NAND2_X1 U417 ( .A1(B[9]), .A2(A[9]), .ZN(n107) );
  NAND2_X1 U418 ( .A1(B[5]), .A2(A[5]), .ZN(n123) );
  NAND2_X1 U419 ( .A1(B[3]), .A2(A[3]), .ZN(n278) );
  NAND2_X1 U420 ( .A1(B[7]), .A2(A[7]), .ZN(n115) );
  NAND2_X1 U421 ( .A1(B[15]), .A2(A[15]), .ZN(n443) );
  NAND2_X1 U422 ( .A1(B[11]), .A2(A[11]), .ZN(n477) );
  OAI21_X1 U423 ( .B1(n231), .B2(n232), .A(n86), .ZN(n199) );
  AND2_X1 U424 ( .A1(A[57]), .A2(B[57]), .ZN(n33) );
  XNOR2_X1 U425 ( .A(n511), .B(n35), .ZN(SUM[53]) );
  OAI21_X1 U426 ( .B1(n34), .B2(net536100), .A(net503746), .ZN(net503770) );
  OAI211_X1 U427 ( .C1(n539), .C2(n329), .A(n332), .B(n331), .ZN(n307) );
  AOI21_X1 U428 ( .B1(net503760), .B2(net503751), .A(n552), .ZN(n168) );
  XNOR2_X1 U429 ( .A(n44), .B(n8), .ZN(SUM[45]) );
  NOR2_X1 U430 ( .A1(n564), .A2(n83), .ZN(n251) );
  AOI21_X1 U431 ( .B1(n236), .B2(n237), .A(n83), .ZN(n231) );
  AOI21_X1 U432 ( .B1(n534), .B2(n160), .A(n547), .ZN(n165) );
  NAND2_X1 U433 ( .A1(n160), .A2(net503708), .ZN(n167) );
  INV_X1 U434 ( .A(n160), .ZN(n546) );
  INV_X1 U435 ( .A(net503753), .ZN(n551) );
  NAND2_X1 U436 ( .A1(net503747), .A2(net503753), .ZN(n35) );
  XNOR2_X1 U437 ( .A(n60), .B(n282), .ZN(SUM[38]) );
  XNOR2_X1 U438 ( .A(n224), .B(n225), .ZN(SUM[47]) );
  AOI21_X1 U439 ( .B1(n226), .B2(n212), .A(n568), .ZN(n224) );
  XNOR2_X1 U440 ( .A(n64), .B(n406), .ZN(SUM[22]) );
  INV_X1 U441 ( .A(n527), .ZN(n136) );
  NOR2_X1 U442 ( .A1(n526), .A2(n527), .ZN(n153) );
  NOR2_X1 U443 ( .A1(B[60]), .A2(A[60]), .ZN(n527) );
  OAI21_X1 U444 ( .B1(n535), .B2(n551), .A(net503747), .ZN(net503760) );
  INV_X1 U445 ( .A(net503770), .ZN(n535) );
  NOR2_X1 U446 ( .A1(B[52]), .A2(A[52]), .ZN(n34) );
  INV_X1 U447 ( .A(n80), .ZN(n572) );
  AND4_X2 U448 ( .A1(n262), .A2(n80), .A3(n263), .A4(n261), .ZN(n76) );
  AND2_X1 U449 ( .A1(B[60]), .A2(A[60]), .ZN(n526) );
  XNOR2_X1 U450 ( .A(n506), .B(n89), .ZN(SUM[28]) );
  NAND2_X1 U451 ( .A1(n65), .A2(n326), .ZN(n357) );
  INV_X1 U452 ( .A(n368), .ZN(n529) );
  INV_X1 U453 ( .A(n219), .ZN(n567) );
  XNOR2_X1 U454 ( .A(n534), .B(n167), .ZN(SUM[58]) );
  NAND2_X1 U455 ( .A1(n404), .A2(n395), .ZN(n403) );
  NAND2_X1 U456 ( .A1(n405), .A2(n398), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n9), .B(n228), .ZN(SUM[46]) );
  NAND2_X1 U458 ( .A1(A[42]), .A2(B[42]), .ZN(n235) );
  AOI21_X1 U459 ( .B1(n159), .B2(net503704), .A(n102), .ZN(n155) );
  NOR2_X1 U460 ( .A1(n521), .A2(n528), .ZN(n148) );
  OR2_X1 U461 ( .A1(n50), .A2(n520), .ZN(n57) );
  XNOR2_X1 U462 ( .A(n520), .B(net503772), .ZN(SUM[52]) );
  OR2_X1 U463 ( .A1(B[37]), .A2(A[37]), .ZN(n262) );
  NOR2_X1 U464 ( .A1(A[37]), .A2(B[37]), .ZN(n266) );
  NAND2_X1 U465 ( .A1(A[37]), .A2(B[37]), .ZN(n269) );
  AND2_X1 U466 ( .A1(B[61]), .A2(A[61]), .ZN(n528) );
  NAND2_X1 U467 ( .A1(n134), .A2(n135), .ZN(n133) );
  NAND2_X1 U468 ( .A1(n514), .A2(n6), .ZN(n194) );
  NAND2_X1 U469 ( .A1(n96), .A2(n87), .ZN(n196) );
  XNOR2_X1 U470 ( .A(n145), .B(n144), .ZN(SUM[62]) );
  NOR2_X1 U471 ( .A1(n300), .A2(n301), .ZN(n299) );
  NAND2_X1 U472 ( .A1(B[63]), .A2(A[63]), .ZN(n130) );
  AND2_X1 U473 ( .A1(n76), .A2(n85), .ZN(n11) );
  NAND2_X1 U474 ( .A1(n76), .A2(n85), .ZN(n259) );
  XNOR2_X1 U475 ( .A(n85), .B(n285), .ZN(SUM[36]) );
  OAI21_X1 U476 ( .B1(n17), .B2(n392), .A(n393), .ZN(n339) );
  XNOR2_X1 U477 ( .A(n254), .B(n255), .ZN(SUM[41]) );
  OAI211_X1 U478 ( .C1(n567), .C2(n208), .A(n209), .B(n210), .ZN(n206) );
  XNOR2_X1 U479 ( .A(n319), .B(n318), .ZN(SUM[33]) );
  NAND2_X1 U480 ( .A1(n294), .A2(n320), .ZN(n319) );
  NAND2_X1 U481 ( .A1(B[56]), .A2(A[56]), .ZN(net503706) );
  XNOR2_X1 U482 ( .A(n250), .B(n251), .ZN(SUM[42]) );
  INV_X1 U483 ( .A(n14), .ZN(n562) );
  AND2_X1 U484 ( .A1(n516), .A2(B[39]), .ZN(n99) );
  OR2_X1 U485 ( .A1(B[39]), .A2(A[39]), .ZN(n80) );
  OAI22_X1 U486 ( .A1(A[39]), .A2(B[39]), .B1(B[38]), .B2(A[38]), .ZN(n38) );
  XNOR2_X1 U487 ( .A(net538671), .B(n48), .ZN(SUM[57]) );
  AOI21_X1 U488 ( .B1(n52), .B2(n53), .A(net534635), .ZN(n51) );
  NAND2_X1 U489 ( .A1(B[54]), .A2(A[54]), .ZN(net503748) );
  OAI21_X1 U490 ( .B1(n22), .B2(n567), .A(n209), .ZN(n9) );
  OAI21_X1 U491 ( .B1(n567), .B2(n22), .A(n209), .ZN(n226) );
  INV_X1 U492 ( .A(n517), .ZN(n563) );
  XNOR2_X1 U493 ( .A(n168), .B(net503756), .ZN(SUM[55]) );
  INV_X1 U494 ( .A(n67), .ZN(n530) );
  XNOR2_X1 U495 ( .A(n391), .B(n67), .ZN(SUM[24]) );
  NAND2_X1 U496 ( .A1(n394), .A2(n393), .ZN(n402) );
  NAND2_X1 U497 ( .A1(n394), .A2(n395), .ZN(n392) );
  AOI21_X1 U498 ( .B1(n229), .B2(n218), .A(n570), .ZN(n22) );
  XNOR2_X1 U499 ( .A(n279), .B(n88), .ZN(SUM[39]) );
  AOI21_X1 U500 ( .B1(n280), .B2(n263), .A(n573), .ZN(n279) );
  AOI21_X1 U501 ( .B1(n260), .B2(n261), .A(n93), .ZN(n95) );
  OAI21_X1 U502 ( .B1(net534627), .B2(n58), .A(net503706), .ZN(net503732) );
  OAI21_X1 U503 ( .B1(n58), .B2(net534627), .A(net503706), .ZN(net538671) );
  INV_X1 U504 ( .A(net503706), .ZN(n550) );
  OAI21_X1 U505 ( .B1(n580), .B2(n537), .A(n399), .ZN(n64) );
  OAI21_X1 U506 ( .B1(n580), .B2(n537), .A(n399), .ZN(n405) );
  NAND2_X1 U507 ( .A1(B[18]), .A2(A[18]), .ZN(n419) );
  OAI21_X1 U508 ( .B1(n531), .B2(n521), .A(n139), .ZN(n144) );
  NOR2_X1 U510 ( .A1(n100), .A2(n102), .ZN(n166) );
  NOR2_X1 U511 ( .A1(n30), .A2(n546), .ZN(n159) );
  NAND2_X1 U512 ( .A1(n130), .A2(n131), .ZN(n128) );
  NAND2_X1 U513 ( .A1(n131), .A2(n143), .ZN(n142) );
  NAND2_X1 U514 ( .A1(n135), .A2(n131), .ZN(n145) );
  NAND2_X1 U515 ( .A1(B[58]), .A2(A[58]), .ZN(net503708) );
  INV_X1 U516 ( .A(n150), .ZN(n531) );
  NOR2_X1 U517 ( .A1(B[59]), .A2(A[59]), .ZN(n100) );
  OAI21_X1 U518 ( .B1(n103), .B2(n245), .A(n246), .ZN(n244) );
  XNOR2_X1 U519 ( .A(n184), .B(n185), .ZN(SUM[51]) );
  AND2_X1 U520 ( .A1(n214), .A2(n213), .ZN(n18) );
  XNOR2_X1 U521 ( .A(n213), .B(n321), .ZN(SUM[32]) );
  NAND2_X1 U522 ( .A1(n213), .A2(n288), .ZN(n287) );
  NAND2_X1 U523 ( .A1(n221), .A2(n213), .ZN(n320) );
  NAND2_X1 U524 ( .A1(B[53]), .A2(A[53]), .ZN(net503747) );
  OAI21_X1 U525 ( .B1(n522), .B2(n527), .A(n140), .ZN(n150) );
  AOI21_X1 U526 ( .B1(n218), .B2(n229), .A(n570), .ZN(n44) );
  XNOR2_X1 U528 ( .A(n230), .B(n508), .ZN(SUM[44]) );
  NAND2_X1 U529 ( .A1(A[43]), .A2(B[43]), .ZN(n234) );
  OAI21_X1 U530 ( .B1(n202), .B2(n75), .A(n199), .ZN(n229) );
  NAND2_X1 U531 ( .A1(n286), .A2(n287), .ZN(n85) );
  NAND2_X1 U532 ( .A1(n286), .A2(n287), .ZN(n260) );
  NAND2_X1 U533 ( .A1(A[35]), .A2(B[35]), .ZN(n297) );
  OR2_X1 U534 ( .A1(A[35]), .A2(B[35]), .ZN(n293) );
  XNOR2_X1 U535 ( .A(n522), .B(n153), .ZN(SUM[60]) );
  NAND2_X1 U536 ( .A1(B[60]), .A2(A[60]), .ZN(n140) );
  XNOR2_X1 U537 ( .A(n42), .B(n409), .ZN(SUM[21]) );
  INV_X1 U538 ( .A(n42), .ZN(n580) );
  NAND2_X1 U539 ( .A1(A[19]), .A2(B[19]), .ZN(n414) );
  AOI21_X1 U540 ( .B1(n205), .B2(n206), .A(n101), .ZN(n195) );
  AOI22_X1 U541 ( .A1(n516), .A2(B[39]), .B1(n571), .B2(n265), .ZN(n14) );
  AND2_X1 U542 ( .A1(n571), .A2(n504), .ZN(n94) );
  NOR2_X1 U543 ( .A1(B[51]), .A2(n501), .ZN(n72) );
  AND2_X1 U544 ( .A1(A[51]), .A2(B[51]), .ZN(n97) );
  OR2_X1 U545 ( .A1(A[51]), .A2(B[51]), .ZN(n176) );
  OAI21_X1 U546 ( .B1(n561), .B2(n95), .A(n525), .ZN(n60) );
  OAI21_X1 U548 ( .B1(n95), .B2(n561), .A(n525), .ZN(n280) );
  XNOR2_X1 U549 ( .A(n148), .B(n531), .ZN(SUM[61]) );
  OAI21_X1 U550 ( .B1(n575), .B2(n204), .A(n76), .ZN(n201) );
  XNOR2_X1 U553 ( .A(n61), .B(n284), .ZN(SUM[37]) );
  INV_X1 U555 ( .A(n41), .ZN(n534) );
  NOR2_X1 U556 ( .A1(n55), .A2(net534635), .ZN(net503756) );
  NOR2_X1 U557 ( .A1(n55), .A2(n553), .ZN(n52) );
  AND2_X1 U559 ( .A1(A[55]), .A2(B[55]), .ZN(net534635) );
  NOR2_X1 U560 ( .A1(A[55]), .A2(B[55]), .ZN(n55) );
  OR2_X1 U561 ( .A1(A[55]), .A2(B[55]), .ZN(net503754) );
  XNOR2_X1 U562 ( .A(n58), .B(n49), .ZN(SUM[56]) );
  NOR2_X1 U563 ( .A1(n550), .A2(net534627), .ZN(n49) );
  AND2_X1 U564 ( .A1(n252), .A2(n253), .ZN(n103) );
  AOI21_X1 U565 ( .B1(n339), .B2(n340), .A(n341), .ZN(n329) );
  AOI21_X1 U566 ( .B1(n4), .B2(n379), .A(n36), .ZN(n74) );
  NAND2_X1 U567 ( .A1(n4), .A2(n379), .ZN(n390) );
  OAI21_X1 U568 ( .B1(n510), .B2(n350), .A(n339), .ZN(n67) );
  OAI21_X1 U569 ( .B1(n510), .B2(n350), .A(n339), .ZN(n4) );
  AOI21_X1 U570 ( .B1(n136), .B2(n137), .A(n138), .ZN(n132) );
  NOR2_X1 U571 ( .A1(B[59]), .A2(A[59]), .ZN(n30) );
  AND2_X1 U572 ( .A1(A[59]), .A2(B[59]), .ZN(n102) );
  AOI21_X1 U573 ( .B1(n186), .B2(n175), .A(n559), .ZN(n184) );
  NAND2_X1 U574 ( .A1(n173), .A2(n513), .ZN(n171) );
  XNOR2_X1 U575 ( .A(n513), .B(n193), .ZN(SUM[48]) );
  XNOR2_X1 U576 ( .A(n186), .B(n188), .ZN(SUM[50]) );
  XNOR2_X1 U577 ( .A(n505), .B(n191), .ZN(SUM[49]) );
  OAI21_X1 U578 ( .B1(n189), .B2(n98), .A(n182), .ZN(n186) );
  AOI21_X1 U579 ( .B1(n172), .B2(n178), .A(n556), .ZN(n189) );
  NAND2_X1 U580 ( .A1(B[45]), .A2(A[45]), .ZN(n209) );
  XNOR2_X1 U581 ( .A(net538470), .B(n169), .ZN(SUM[54]) );
  OAI21_X1 U582 ( .B1(n551), .B2(n535), .A(net503747), .ZN(net538470) );
  NOR2_X1 U583 ( .A1(n509), .A2(net534627), .ZN(net503696) );
  OAI211_X1 U584 ( .C1(n509), .C2(net503706), .A(n549), .B(net503708), .ZN(
        net503704) );
  INV_X1 U585 ( .A(net534734), .ZN(n548) );
  OR2_X1 U586 ( .A1(n33), .A2(net534734), .ZN(n48) );
  NOR2_X1 U587 ( .A1(n100), .A2(n546), .ZN(n157) );
  XNOR2_X1 U588 ( .A(n166), .B(n165), .ZN(SUM[59]) );
endmodule


module RCA_NBIT64_7 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_7_DW01_add_6 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_6_DW01_add_8 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net489131, net489130, net489114, net489101, net489093, net489091,
         net489134, net489125, net489099, net489092, net489122, net489120,
         net489106, net489105, net537531, net489126, net489103, net489128, n2,
         n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n20,
         n22, n25, n28, n29, n30, n31, n36, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n50, n51, n52, n53, n54, n56, n58, n59, n60, n61, n62, n63,
         n64, n65, n69, n70, n71, n72, n73, n74, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n97,
         n98, n99, n100, n102, n103, n104, n105, n106, n107, n110, n111, n113,
         n114, n115, n117, n119, n121, n122, n123, n124, n125, n126, n127,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n144, n146, n147, n148, n150, n151, n152, n153,
         n154, n155, n156, n157, n160, n161, n162, n163, n164, n165, n166,
         n168, n169, n170, n171, n172, n173, n174, n175, n177, n179, n180,
         n181, n182, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n200, n201, n202, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n220,
         n221, n222, n223, n224, n226, n227, n228, n229, n230, n231, n233,
         n234, n235, n237, n238, n239, n240, n242, n243, n246, n247, n248,
         n249, n252, n254, n255, n256, n257, n258, n259, n263, n264, n265,
         n268, n271, n272, n273, n274, n275, n277, n278, n283, n284, n285,
         n286, n287, n288, n289, n291, n292, n293, n295, n296, n297, n298,
         n299, n303, n304, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n318, n319, n320, n321, n323, n324, n325, n326, n329, n330,
         n331, n332, n334, n335, n336, n337, n338, n339, n340, n342, n343,
         n344, n347, n348, n349, n350, n352, n353, n354, n355, n357, n358,
         n359, n360, n361, n362, n363, n365, n367, n368, n371, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n417, n418, n419, n420, n421, n422,
         n424, n425, n426, n427, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n447, n448,
         n450, n451, n455, n456, n457, n458, n459, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n474, n475, n477,
         n478, n479, n480, n481, n482, n484, n486, n487, n488, n489, n490,
         n493, n494, n495, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n529,
         n530, n531, n532, n534, n536, n537, n538, n539, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660;

  NAND3_X1 U6 ( .A1(n227), .A2(n226), .A3(n3), .ZN(n193) );
  NAND3_X1 U17 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n9) );
  OR2_X2 U26 ( .A1(A[34]), .A2(B[34]), .ZN(n46) );
  NAND3_X1 U44 ( .A1(n216), .A2(n220), .A3(n284), .ZN(n252) );
  OR2_X2 U113 ( .A1(A[54]), .A2(B[54]), .ZN(n140) );
  OR2_X2 U360 ( .A1(B[44]), .A2(A[44]), .ZN(n214) );
  OR2_X2 U362 ( .A1(A[45]), .A2(B[45]), .ZN(n213) );
  OR2_X2 U363 ( .A1(B[49]), .A2(A[49]), .ZN(n164) );
  OR2_X2 U364 ( .A1(B[48]), .A2(A[48]), .ZN(n174) );
  OR2_X2 U367 ( .A1(B[29]), .A2(A[29]), .ZN(n375) );
  OR2_X2 U376 ( .A1(B[40]), .A2(A[40]), .ZN(n265) );
  NAND3_X1 U527 ( .A1(n152), .A2(n148), .A3(n153), .ZN(n151) );
  NAND3_X1 U528 ( .A1(n154), .A2(n140), .A3(n135), .ZN(n153) );
  NAND3_X1 U533 ( .A1(n162), .A2(n177), .A3(n163), .ZN(n175) );
  NAND3_X1 U534 ( .A1(A[48]), .A2(B[48]), .A3(n164), .ZN(n177) );
  NAND3_X1 U535 ( .A1(n47), .A2(n5), .A3(n174), .ZN(n180) );
  NAND3_X1 U538 ( .A1(n264), .A2(n213), .A3(n214), .ZN(n208) );
  NAND3_X1 U550 ( .A1(n248), .A2(n247), .A3(n201), .ZN(n238) );
  NAND3_X1 U553 ( .A1(n226), .A2(n252), .A3(n214), .ZN(n247) );
  NAND3_X1 U556 ( .A1(n256), .A2(n255), .A3(n254), .ZN(n206) );
  NAND3_X1 U557 ( .A1(n259), .A2(n263), .A3(n618), .ZN(n255) );
  NAND3_X1 U566 ( .A1(n291), .A2(n220), .A3(n284), .ZN(n289) );
  NAND3_X1 U574 ( .A1(n293), .A2(n554), .A3(n560), .ZN(n216) );
  NAND3_X1 U575 ( .A1(n304), .A2(n303), .A3(n621), .ZN(n293) );
  NAND3_X1 U580 ( .A1(n330), .A2(n329), .A3(n46), .ZN(n342) );
  NAND3_X1 U584 ( .A1(n548), .A2(n329), .A3(n324), .ZN(n350) );
  NAND3_X1 U588 ( .A1(n550), .A2(n376), .A3(n377), .ZN(n353) );
  NAND3_X1 U594 ( .A1(n392), .A2(n390), .A3(n391), .ZN(n396) );
  NAND3_X1 U595 ( .A1(n380), .A2(n360), .A3(n361), .ZN(n391) );
  NAND3_X1 U596 ( .A1(n380), .A2(n403), .A3(n382), .ZN(n392) );
  NAND3_X1 U599 ( .A1(n407), .A2(n408), .A3(n409), .ZN(n406) );
  NAND3_X1 U624 ( .A1(n517), .A2(n518), .A3(n519), .ZN(n516) );
  NAND3_X1 U625 ( .A1(n520), .A2(n80), .A3(n521), .ZN(n517) );
  OR2_X2 U8 ( .A1(A[46]), .A2(B[46]), .ZN(n210) );
  OR2_X2 U18 ( .A1(A[58]), .A2(B[58]), .ZN(net489106) );
  OR2_X2 U378 ( .A1(B[36]), .A2(A[36]), .ZN(n228) );
  OR2_X2 U2 ( .A1(A[43]), .A2(B[43]), .ZN(n264) );
  CLKBUF_X1 U3 ( .A(A[43]), .Z(n542) );
  OR2_X1 U4 ( .A1(n44), .A2(n609), .ZN(n190) );
  OR2_X1 U5 ( .A1(B[53]), .A2(A[53]), .ZN(n138) );
  OR2_X1 U7 ( .A1(B[52]), .A2(A[52]), .ZN(n137) );
  AND2_X1 U9 ( .A1(n534), .A2(n467), .ZN(SUM[0]) );
  OR2_X1 U10 ( .A1(B[56]), .A2(A[56]), .ZN(net489099) );
  CLKBUF_X1 U11 ( .A(A[35]), .Z(n543) );
  AND2_X1 U12 ( .A1(A[41]), .A2(B[41]), .ZN(n544) );
  AND2_X1 U13 ( .A1(net489092), .A2(n556), .ZN(n545) );
  AND2_X1 U14 ( .A1(n136), .A2(n135), .ZN(n546) );
  NOR2_X1 U15 ( .A1(n209), .A2(n208), .ZN(n547) );
  BUF_X2 U16 ( .A(n326), .Z(n548) );
  OAI221_X1 U19 ( .B1(n325), .B2(n60), .C1(n629), .C2(n625), .A(n222), .ZN(
        n549) );
  NAND2_X1 U20 ( .A1(n656), .A2(n581), .ZN(n550) );
  NOR2_X1 U21 ( .A1(B[53]), .A2(A[53]), .ZN(n551) );
  OR2_X2 U22 ( .A1(A[57]), .A2(B[57]), .ZN(net489128) );
  OR2_X2 U23 ( .A1(B[37]), .A2(A[37]), .ZN(n229) );
  NAND2_X1 U24 ( .A1(n259), .A2(n544), .ZN(n254) );
  AND3_X2 U25 ( .A1(n212), .A2(n7), .A3(n14), .ZN(n226) );
  NAND3_X1 U27 ( .A1(n248), .A2(n247), .A3(n201), .ZN(n552) );
  AOI21_X1 U28 ( .B1(n141), .B2(n142), .A(n599), .ZN(n553) );
  OR2_X1 U29 ( .A1(A[39]), .A2(B[39]), .ZN(n554) );
  OR2_X1 U30 ( .A1(A[39]), .A2(B[39]), .ZN(n231) );
  NOR2_X1 U31 ( .A1(B[33]), .A2(A[33]), .ZN(n555) );
  OR2_X1 U32 ( .A1(B[33]), .A2(A[33]), .ZN(n330) );
  NAND2_X1 U33 ( .A1(n330), .A2(n336), .ZN(n349) );
  NAND2_X1 U34 ( .A1(n553), .A2(n133), .ZN(n556) );
  AND2_X1 U35 ( .A1(n164), .A2(n174), .ZN(n557) );
  AND3_X1 U36 ( .A1(n172), .A2(n559), .A3(n557), .ZN(n171) );
  XNOR2_X1 U37 ( .A(n268), .B(n558), .ZN(SUM[43]) );
  NOR2_X1 U38 ( .A1(n77), .A2(n561), .ZN(n558) );
  OAI21_X2 U39 ( .B1(n636), .B2(n368), .A(n367), .ZN(n403) );
  OR2_X2 U40 ( .A1(B[22]), .A2(A[22]), .ZN(n435) );
  NAND2_X1 U41 ( .A1(n134), .A2(n546), .ZN(n133) );
  OR2_X1 U42 ( .A1(B[50]), .A2(A[50]), .ZN(n559) );
  OR2_X1 U43 ( .A1(A[50]), .A2(B[50]), .ZN(n173) );
  NAND2_X1 U45 ( .A1(A[45]), .A2(B[45]), .ZN(n240) );
  OR2_X1 U46 ( .A1(B[42]), .A2(A[42]), .ZN(n7) );
  OR2_X1 U47 ( .A1(B[41]), .A2(A[41]), .ZN(n263) );
  AND2_X1 U48 ( .A1(n62), .A2(n63), .ZN(n560) );
  INV_X1 U49 ( .A(n264), .ZN(n561) );
  AND2_X1 U50 ( .A1(n148), .A2(n140), .ZN(n157) );
  NAND2_X1 U51 ( .A1(n565), .A2(n169), .ZN(n562) );
  AND2_X1 U52 ( .A1(n562), .A2(n563), .ZN(n166) );
  OR2_X1 U53 ( .A1(n564), .A2(n137), .ZN(n563) );
  INV_X1 U54 ( .A(n146), .ZN(n564) );
  AND2_X1 U55 ( .A1(n161), .A2(n146), .ZN(n565) );
  INV_X1 U56 ( .A(n620), .ZN(n566) );
  NAND2_X1 U57 ( .A1(n126), .A2(n545), .ZN(net489091) );
  XOR2_X1 U58 ( .A(n22), .B(n567), .Z(SUM[39]) );
  NAND2_X1 U59 ( .A1(n554), .A2(n220), .ZN(n567) );
  XNOR2_X1 U60 ( .A(n179), .B(n568), .ZN(SUM[51]) );
  NAND2_X1 U61 ( .A1(n160), .A2(n59), .ZN(n568) );
  INV_X1 U62 ( .A(n450), .ZN(n636) );
  NAND2_X1 U63 ( .A1(n331), .A2(n332), .ZN(n221) );
  NOR2_X1 U64 ( .A1(n612), .A2(n607), .ZN(n237) );
  INV_X1 U65 ( .A(n293), .ZN(n603) );
  NOR2_X1 U66 ( .A1(n619), .A2(n624), .ZN(n278) );
  NOR2_X1 U67 ( .A1(n615), .A2(n619), .ZN(n288) );
  INV_X1 U68 ( .A(A[26]), .ZN(n578) );
  INV_X1 U69 ( .A(n275), .ZN(n615) );
  INV_X1 U70 ( .A(n447), .ZN(n634) );
  INV_X1 U71 ( .A(n223), .ZN(n606) );
  INV_X1 U72 ( .A(n123), .ZN(n573) );
  INV_X1 U73 ( .A(n284), .ZN(n575) );
  OAI21_X1 U74 ( .B1(n658), .B2(n502), .A(n499), .ZN(n83) );
  OAI21_X1 U75 ( .B1(n642), .B2(n383), .A(n637), .ZN(n450) );
  INV_X1 U76 ( .A(n365), .ZN(n637) );
  AOI21_X1 U77 ( .B1(n498), .B2(n499), .A(n500), .ZN(n495) );
  NAND2_X1 U78 ( .A1(n650), .A2(n501), .ZN(n498) );
  INV_X1 U79 ( .A(n502), .ZN(n650) );
  NOR2_X1 U80 ( .A1(n383), .A2(n368), .ZN(n381) );
  NAND2_X1 U81 ( .A1(n514), .A2(n497), .ZN(n512) );
  NAND2_X1 U82 ( .A1(n646), .A2(n83), .ZN(n514) );
  INV_X1 U83 ( .A(n500), .ZN(n646) );
  INV_X1 U84 ( .A(n368), .ZN(n632) );
  INV_X1 U85 ( .A(n501), .ZN(n658) );
  INV_X1 U86 ( .A(n376), .ZN(n642) );
  NOR2_X1 U87 ( .A1(n100), .A2(n590), .ZN(SUM[64]) );
  INV_X1 U88 ( .A(n497), .ZN(n647) );
  NOR2_X1 U89 ( .A1(n610), .A2(n609), .ZN(n65) );
  AOI21_X1 U90 ( .B1(n237), .B2(n552), .A(n239), .ZN(n235) );
  INV_X1 U91 ( .A(n191), .ZN(n610) );
  XOR2_X1 U92 ( .A(n19), .B(n569), .Z(SUM[32]) );
  NAND2_X1 U93 ( .A1(n334), .A2(n329), .ZN(n569) );
  NOR2_X1 U94 ( .A1(n617), .A2(n615), .ZN(n296) );
  XNOR2_X1 U95 ( .A(n349), .B(n570), .ZN(SUM[33]) );
  NAND2_X1 U96 ( .A1(n350), .A2(n334), .ZN(n570) );
  NAND2_X1 U97 ( .A1(n265), .A2(n285), .ZN(n297) );
  NAND2_X1 U98 ( .A1(n373), .A2(n326), .ZN(n2) );
  AND4_X1 U99 ( .A1(n389), .A2(n390), .A3(n391), .A4(n392), .ZN(n11) );
  NAND2_X1 U100 ( .A1(n318), .A2(n230), .ZN(n320) );
  NAND2_X1 U101 ( .A1(n8), .A2(n144), .ZN(n150) );
  NAND2_X1 U102 ( .A1(n413), .A2(n411), .ZN(n427) );
  XOR2_X1 U103 ( .A(n170), .B(n571), .Z(SUM[48]) );
  AND2_X1 U104 ( .A1(n174), .A2(n184), .ZN(n571) );
  NOR2_X1 U105 ( .A1(n627), .A2(n628), .ZN(n344) );
  NOR2_X1 U106 ( .A1(n347), .A2(n626), .ZN(n343) );
  INV_X1 U107 ( .A(n335), .ZN(n627) );
  OAI21_X1 U108 ( .B1(n605), .B2(n574), .A(n307), .ZN(n52) );
  INV_X1 U109 ( .A(n228), .ZN(n605) );
  XNOR2_X1 U110 ( .A(n238), .B(n246), .ZN(SUM[45]) );
  NAND2_X1 U111 ( .A1(n213), .A2(n240), .ZN(n246) );
  OAI211_X1 U112 ( .C1(n325), .C2(n60), .A(n222), .B(n221), .ZN(n299) );
  NOR2_X1 U114 ( .A1(n608), .A2(n607), .ZN(n243) );
  AOI21_X1 U115 ( .B1(n213), .B2(n552), .A(n611), .ZN(n242) );
  INV_X1 U116 ( .A(n202), .ZN(n608) );
  INV_X1 U117 ( .A(n411), .ZN(n577) );
  XNOR2_X1 U118 ( .A(n136), .B(n168), .ZN(SUM[52]) );
  NAND2_X1 U119 ( .A1(n146), .A2(n137), .ZN(n168) );
  AOI21_X1 U120 ( .B1(n113), .B2(n115), .A(n591), .ZN(n114) );
  INV_X1 U121 ( .A(n107), .ZN(n591) );
  XNOR2_X1 U122 ( .A(n195), .B(n196), .ZN(SUM[49]) );
  NOR2_X1 U123 ( .A1(n72), .A2(n587), .ZN(n196) );
  AOI21_X1 U124 ( .B1(n47), .B2(n174), .A(n600), .ZN(n195) );
  INV_X1 U125 ( .A(n164), .ZN(n587) );
  NAND4_X1 U126 ( .A1(n193), .A2(n36), .A3(n190), .A4(n191), .ZN(n47) );
  NAND2_X1 U127 ( .A1(n207), .A2(n53), .ZN(n36) );
  INV_X1 U128 ( .A(net489106), .ZN(n595) );
  XNOR2_X1 U129 ( .A(n402), .B(n396), .ZN(SUM[29]) );
  NAND2_X1 U130 ( .A1(n375), .A2(n389), .ZN(n402) );
  XNOR2_X1 U131 ( .A(n299), .B(n323), .ZN(SUM[36]) );
  NAND2_X1 U132 ( .A1(n228), .A2(n307), .ZN(n323) );
  XNOR2_X1 U133 ( .A(n404), .B(n45), .ZN(SUM[28]) );
  NOR2_X1 U134 ( .A1(n582), .A2(n583), .ZN(n45) );
  INV_X1 U135 ( .A(n380), .ZN(n583) );
  XNOR2_X1 U136 ( .A(n444), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U137 ( .A1(n435), .A2(n433), .ZN(n444) );
  OAI21_X1 U138 ( .B1(n634), .B2(n633), .A(n437), .ZN(n16) );
  XNOR2_X1 U139 ( .A(n425), .B(n424), .ZN(SUM[25]) );
  NAND2_X1 U140 ( .A1(n426), .A2(n411), .ZN(n424) );
  AND2_X1 U141 ( .A1(n606), .A2(n224), .ZN(n3) );
  AND2_X1 U142 ( .A1(n30), .A2(n41), .ZN(n227) );
  XNOR2_X1 U143 ( .A(n441), .B(n440), .ZN(SUM[23]) );
  NAND2_X1 U144 ( .A1(n433), .A2(n442), .ZN(n441) );
  NAND2_X1 U145 ( .A1(n443), .A2(n435), .ZN(n442) );
  OAI21_X1 U146 ( .B1(n430), .B2(n429), .A(n431), .ZN(n367) );
  NAND2_X1 U147 ( .A1(n437), .A2(n438), .ZN(n436) );
  AND2_X1 U148 ( .A1(n285), .A2(n286), .ZN(n272) );
  NAND2_X1 U149 ( .A1(n275), .A2(n7), .ZN(n274) );
  AOI21_X1 U150 ( .B1(n221), .B2(n222), .A(n223), .ZN(n218) );
  OAI211_X1 U151 ( .C1(n70), .C2(n584), .A(n161), .B(n160), .ZN(n154) );
  AND3_X1 U152 ( .A1(n162), .A2(n177), .A3(n163), .ZN(n70) );
  AOI21_X1 U153 ( .B1(n233), .B2(n334), .A(n348), .ZN(n347) );
  NAND4_X1 U154 ( .A1(n298), .A2(n231), .A3(n228), .A4(n299), .ZN(n284) );
  AOI21_X1 U155 ( .B1(n621), .B2(n655), .A(n620), .ZN(n298) );
  AND2_X1 U156 ( .A1(n329), .A2(n330), .ZN(n56) );
  NAND2_X1 U157 ( .A1(n656), .A2(n581), .ZN(n374) );
  OAI211_X1 U158 ( .C1(n146), .C2(n551), .A(n147), .B(n148), .ZN(n142) );
  AOI21_X1 U159 ( .B1(n215), .B2(n216), .A(n217), .ZN(n205) );
  NOR2_X1 U160 ( .A1(n218), .A2(n623), .ZN(n215) );
  NAND4_X1 U161 ( .A1(n263), .A2(n264), .A3(n265), .A4(n7), .ZN(n217) );
  XNOR2_X1 U162 ( .A(n39), .B(n40), .ZN(SUM[44]) );
  OR2_X1 U163 ( .A1(n613), .A2(n614), .ZN(n40) );
  NAND2_X1 U164 ( .A1(n42), .A2(n43), .ZN(n39) );
  INV_X1 U165 ( .A(n201), .ZN(n613) );
  XNOR2_X1 U166 ( .A(n418), .B(n417), .ZN(SUM[27]) );
  NAND2_X1 U167 ( .A1(n360), .A2(n421), .ZN(n417) );
  NAND2_X1 U168 ( .A1(n419), .A2(n412), .ZN(n418) );
  OAI21_X1 U169 ( .B1(n551), .B2(n146), .A(n147), .ZN(n155) );
  OAI21_X1 U170 ( .B1(n635), .B2(n636), .A(n438), .ZN(n447) );
  INV_X1 U171 ( .A(n439), .ZN(n635) );
  OAI21_X1 U172 ( .B1(n628), .B2(n336), .A(n335), .ZN(n340) );
  OAI21_X1 U173 ( .B1(n607), .B2(n240), .A(n202), .ZN(n239) );
  OAI21_X1 U174 ( .B1(n634), .B2(n633), .A(n437), .ZN(n443) );
  NAND2_X1 U175 ( .A1(n362), .A2(n363), .ZN(n382) );
  NAND2_X1 U176 ( .A1(n405), .A2(n406), .ZN(n361) );
  AND2_X1 U177 ( .A1(n421), .A2(n412), .ZN(n405) );
  NAND2_X1 U178 ( .A1(n410), .A2(n411), .ZN(n408) );
  XNOR2_X1 U179 ( .A(n448), .B(n447), .ZN(SUM[21]) );
  AOI21_X1 U180 ( .B1(n292), .B2(n283), .A(n618), .ZN(n291) );
  NOR2_X1 U181 ( .A1(n624), .A2(n603), .ZN(n292) );
  INV_X1 U182 ( .A(n210), .ZN(n607) );
  OAI21_X1 U183 ( .B1(n602), .B2(n603), .A(n220), .ZN(n277) );
  INV_X1 U184 ( .A(n283), .ZN(n602) );
  NAND2_X1 U185 ( .A1(n657), .A2(n578), .ZN(n409) );
  NAND2_X1 U186 ( .A1(n621), .A2(n655), .ZN(n230) );
  AND2_X1 U187 ( .A1(n337), .A2(n222), .ZN(n50) );
  NOR2_X1 U188 ( .A1(n339), .A2(n340), .ZN(n338) );
  NAND2_X1 U189 ( .A1(n654), .A2(n616), .ZN(n275) );
  XNOR2_X1 U190 ( .A(n393), .B(n394), .ZN(SUM[30]) );
  NAND2_X1 U191 ( .A1(n374), .A2(n386), .ZN(n393) );
  NAND2_X1 U192 ( .A1(n395), .A2(n389), .ZN(n394) );
  NAND2_X1 U193 ( .A1(n375), .A2(n396), .ZN(n395) );
  AND2_X1 U194 ( .A1(n263), .A2(n265), .ZN(n14) );
  NAND2_X1 U195 ( .A1(n200), .A2(n210), .ZN(n44) );
  OAI211_X1 U196 ( .C1(n612), .C2(n201), .A(n240), .B(n202), .ZN(n200) );
  AND2_X1 U197 ( .A1(n337), .A2(n46), .ZN(n331) );
  NOR2_X1 U198 ( .A1(n182), .A2(n586), .ZN(n181) );
  INV_X1 U199 ( .A(n162), .ZN(n586) );
  NOR2_X1 U200 ( .A1(n58), .A2(n185), .ZN(n182) );
  AND2_X1 U201 ( .A1(n163), .A2(n184), .ZN(n58) );
  NAND2_X1 U202 ( .A1(n329), .A2(n330), .ZN(n348) );
  NOR2_X1 U203 ( .A1(n593), .A2(n598), .ZN(net489092) );
  INV_X1 U204 ( .A(net489099), .ZN(n598) );
  INV_X1 U205 ( .A(net489128), .ZN(n593) );
  INV_X1 U206 ( .A(n285), .ZN(n618) );
  INV_X1 U207 ( .A(n265), .ZN(n619) );
  INV_X1 U208 ( .A(n231), .ZN(n624) );
  XNOR2_X1 U209 ( .A(n31), .B(n422), .ZN(SUM[26]) );
  NAND2_X1 U210 ( .A1(n412), .A2(n409), .ZN(n422) );
  INV_X1 U211 ( .A(n46), .ZN(n628) );
  INV_X1 U212 ( .A(n213), .ZN(n612) );
  OAI221_X1 U213 ( .B1(n325), .B2(n60), .C1(n629), .C2(n625), .A(n222), .ZN(
        n28) );
  INV_X1 U214 ( .A(n331), .ZN(n629) );
  INV_X1 U215 ( .A(n332), .ZN(n625) );
  NAND2_X1 U216 ( .A1(n384), .A2(n550), .ZN(n352) );
  NAND2_X1 U217 ( .A1(n389), .A2(n386), .ZN(n384) );
  NAND2_X1 U218 ( .A1(n547), .A2(n53), .ZN(n192) );
  INV_X1 U219 ( .A(n286), .ZN(n617) );
  NAND2_X1 U220 ( .A1(n580), .A2(n357), .ZN(n355) );
  OAI21_X1 U221 ( .B1(n358), .B2(n69), .A(n359), .ZN(n357) );
  INV_X1 U222 ( .A(n25), .ZN(n580) );
  AOI21_X1 U223 ( .B1(n632), .B2(n365), .A(n631), .ZN(n358) );
  INV_X1 U224 ( .A(n390), .ZN(n582) );
  NAND2_X1 U225 ( .A1(n206), .A2(n264), .ZN(n43) );
  NAND2_X1 U226 ( .A1(n657), .A2(n578), .ZN(n414) );
  NAND2_X1 U227 ( .A1(n360), .A2(n361), .ZN(n359) );
  INV_X1 U228 ( .A(n30), .ZN(n609) );
  NAND2_X1 U229 ( .A1(n189), .A2(n174), .ZN(n188) );
  INV_X1 U230 ( .A(n240), .ZN(n611) );
  INV_X1 U231 ( .A(n220), .ZN(n623) );
  INV_X1 U232 ( .A(n336), .ZN(n626) );
  NAND2_X1 U233 ( .A1(n375), .A2(n374), .ZN(n388) );
  INV_X1 U234 ( .A(n307), .ZN(n604) );
  INV_X1 U235 ( .A(n184), .ZN(n600) );
  AND2_X1 U236 ( .A1(n362), .A2(n363), .ZN(n69) );
  AND2_X1 U237 ( .A1(n13), .A2(n210), .ZN(n41) );
  AND3_X1 U238 ( .A1(n46), .A2(n214), .A3(n213), .ZN(n13) );
  INV_X1 U239 ( .A(n214), .ZN(n614) );
  NAND2_X1 U240 ( .A1(n61), .A2(n324), .ZN(n60) );
  AND2_X1 U241 ( .A1(n46), .A2(n548), .ZN(n61) );
  INV_X1 U242 ( .A(n318), .ZN(n622) );
  AND2_X1 U243 ( .A1(n8), .A2(n140), .ZN(n134) );
  AND2_X1 U244 ( .A1(n360), .A2(n361), .ZN(n12) );
  XNOR2_X1 U245 ( .A(n503), .B(n504), .ZN(SUM[15]) );
  NAND2_X1 U246 ( .A1(n505), .A2(n488), .ZN(n504) );
  NAND2_X1 U247 ( .A1(n484), .A2(n490), .ZN(n503) );
  NAND2_X1 U248 ( .A1(n489), .A2(n506), .ZN(n505) );
  XNOR2_X1 U249 ( .A(n451), .B(n450), .ZN(SUM[20]) );
  NAND2_X1 U250 ( .A1(n439), .A2(n438), .ZN(n451) );
  XNOR2_X1 U251 ( .A(n475), .B(n474), .ZN(SUM[17]) );
  NAND2_X1 U252 ( .A1(n465), .A2(n462), .ZN(n475) );
  XNOR2_X1 U253 ( .A(n468), .B(n469), .ZN(SUM[19]) );
  NAND2_X1 U254 ( .A1(n463), .A2(n470), .ZN(n469) );
  NAND2_X1 U255 ( .A1(n458), .A2(n456), .ZN(n468) );
  NAND2_X1 U256 ( .A1(n457), .A2(n471), .ZN(n470) );
  XNOR2_X1 U257 ( .A(n472), .B(n471), .ZN(SUM[18]) );
  NAND2_X1 U258 ( .A1(n457), .A2(n463), .ZN(n472) );
  XNOR2_X1 U259 ( .A(n507), .B(n506), .ZN(SUM[14]) );
  NAND2_X1 U260 ( .A1(n489), .A2(n488), .ZN(n507) );
  XNOR2_X1 U261 ( .A(n510), .B(n509), .ZN(SUM[13]) );
  NAND2_X1 U262 ( .A1(n494), .A2(n487), .ZN(n510) );
  XNOR2_X1 U263 ( .A(n477), .B(n376), .ZN(SUM[16]) );
  NAND2_X1 U264 ( .A1(n464), .A2(n461), .ZN(n477) );
  XNOR2_X1 U265 ( .A(n86), .B(n87), .ZN(SUM[7]) );
  NAND2_X1 U266 ( .A1(n90), .A2(n91), .ZN(n86) );
  NAND2_X1 U267 ( .A1(n88), .A2(n89), .ZN(n87) );
  NAND2_X1 U268 ( .A1(n92), .A2(n93), .ZN(n91) );
  XNOR2_X1 U269 ( .A(n308), .B(n309), .ZN(SUM[3]) );
  NAND2_X1 U270 ( .A1(n312), .A2(n313), .ZN(n308) );
  NAND2_X1 U271 ( .A1(n310), .A2(n311), .ZN(n309) );
  NAND2_X1 U272 ( .A1(n314), .A2(n315), .ZN(n313) );
  XNOR2_X1 U273 ( .A(n522), .B(n523), .ZN(SUM[11]) );
  NAND2_X1 U274 ( .A1(n518), .A2(n524), .ZN(n523) );
  NAND2_X1 U275 ( .A1(n519), .A2(n515), .ZN(n522) );
  NAND2_X1 U276 ( .A1(n521), .A2(n525), .ZN(n524) );
  XNOR2_X1 U277 ( .A(n466), .B(n660), .ZN(SUM[1]) );
  NAND2_X1 U278 ( .A1(n400), .A2(n399), .ZN(n466) );
  XNOR2_X1 U279 ( .A(n513), .B(n512), .ZN(SUM[12]) );
  NAND2_X1 U280 ( .A1(n493), .A2(n486), .ZN(n513) );
  XNOR2_X1 U281 ( .A(n82), .B(n83), .ZN(SUM[8]) );
  NAND2_X1 U282 ( .A1(n84), .A2(n85), .ZN(n82) );
  XNOR2_X1 U283 ( .A(n78), .B(n79), .ZN(SUM[9]) );
  NAND2_X1 U284 ( .A1(n80), .A2(n81), .ZN(n78) );
  XNOR2_X1 U285 ( .A(n127), .B(n99), .ZN(SUM[5]) );
  NAND2_X1 U286 ( .A1(n98), .A2(n97), .ZN(n127) );
  XNOR2_X1 U287 ( .A(n94), .B(n92), .ZN(SUM[6]) );
  NAND2_X1 U288 ( .A1(n93), .A2(n90), .ZN(n94) );
  XNOR2_X1 U289 ( .A(n526), .B(n525), .ZN(SUM[10]) );
  NAND2_X1 U290 ( .A1(n521), .A2(n518), .ZN(n526) );
  XNOR2_X1 U291 ( .A(n397), .B(n314), .ZN(SUM[2]) );
  NAND2_X1 U292 ( .A1(n315), .A2(n312), .ZN(n397) );
  XNOR2_X1 U293 ( .A(n194), .B(n501), .ZN(SUM[4]) );
  NAND2_X1 U294 ( .A1(n130), .A2(n129), .ZN(n194) );
  OAI21_X1 U295 ( .B1(n536), .B2(n537), .A(n311), .ZN(n501) );
  NAND2_X1 U296 ( .A1(n315), .A2(n310), .ZN(n537) );
  NOR2_X1 U297 ( .A1(n538), .A2(n539), .ZN(n536) );
  NAND2_X1 U298 ( .A1(n312), .A2(n399), .ZN(n539) );
  OAI21_X1 U299 ( .B1(n478), .B2(n479), .A(n480), .ZN(n376) );
  NOR2_X1 U300 ( .A1(n495), .A2(n647), .ZN(n478) );
  NAND4_X1 U301 ( .A1(n493), .A2(n494), .A3(n489), .A4(n490), .ZN(n479) );
  AOI21_X1 U302 ( .B1(n481), .B2(n482), .A(n643), .ZN(n480) );
  OAI21_X1 U303 ( .B1(n649), .B2(n648), .A(n81), .ZN(n525) );
  INV_X1 U304 ( .A(n79), .ZN(n649) );
  INV_X1 U305 ( .A(n80), .ZN(n648) );
  OAI21_X1 U306 ( .B1(n645), .B2(n644), .A(n487), .ZN(n506) );
  INV_X1 U307 ( .A(n509), .ZN(n645) );
  OAI21_X1 U308 ( .B1(n640), .B2(n639), .A(n462), .ZN(n471) );
  INV_X1 U309 ( .A(n474), .ZN(n640) );
  OAI21_X1 U310 ( .B1(n642), .B2(n641), .A(n461), .ZN(n474) );
  INV_X1 U311 ( .A(n464), .ZN(n641) );
  OAI21_X1 U312 ( .B1(n653), .B2(n658), .A(n129), .ZN(n99) );
  INV_X1 U313 ( .A(n130), .ZN(n653) );
  OAI21_X1 U314 ( .B1(n652), .B2(n651), .A(n97), .ZN(n92) );
  INV_X1 U315 ( .A(n99), .ZN(n652) );
  INV_X1 U316 ( .A(n98), .ZN(n651) );
  OAI21_X1 U317 ( .B1(n638), .B2(n455), .A(n456), .ZN(n365) );
  INV_X1 U318 ( .A(n459), .ZN(n638) );
  NAND2_X1 U319 ( .A1(n457), .A2(n458), .ZN(n455) );
  OAI211_X1 U320 ( .C1(n639), .C2(n461), .A(n462), .B(n463), .ZN(n459) );
  OAI21_X1 U321 ( .B1(n530), .B2(n531), .A(n88), .ZN(n499) );
  NAND2_X1 U322 ( .A1(n89), .A2(n90), .ZN(n531) );
  NOR2_X1 U323 ( .A1(n15), .A2(n532), .ZN(n530) );
  AND2_X1 U324 ( .A1(n97), .A2(n129), .ZN(n15) );
  NAND4_X1 U325 ( .A1(n464), .A2(n465), .A3(n457), .A4(n458), .ZN(n383) );
  NAND4_X1 U326 ( .A1(n130), .A2(n98), .A3(n93), .A4(n88), .ZN(n502) );
  NAND4_X1 U327 ( .A1(n80), .A2(n84), .A3(n521), .A4(n515), .ZN(n500) );
  AOI21_X1 U328 ( .B1(n103), .B2(n104), .A(n105), .ZN(n100) );
  NAND2_X1 U329 ( .A1(n106), .A2(n107), .ZN(n105) );
  NOR2_X1 U330 ( .A1(n592), .A2(n71), .ZN(n103) );
  OAI211_X1 U331 ( .C1(n644), .C2(n486), .A(n487), .B(n488), .ZN(n482) );
  NOR2_X1 U332 ( .A1(n378), .A2(n379), .ZN(n377) );
  NAND2_X1 U333 ( .A1(n381), .A2(n382), .ZN(n378) );
  NAND2_X1 U334 ( .A1(n380), .A2(n375), .ZN(n379) );
  NOR2_X1 U335 ( .A1(n659), .A2(n467), .ZN(n538) );
  INV_X1 U336 ( .A(n400), .ZN(n659) );
  NAND2_X1 U337 ( .A1(n529), .A2(n85), .ZN(n79) );
  NAND2_X1 U338 ( .A1(n83), .A2(n84), .ZN(n529) );
  NAND2_X1 U339 ( .A1(n511), .A2(n486), .ZN(n509) );
  NAND2_X1 U340 ( .A1(n512), .A2(n493), .ZN(n511) );
  NAND2_X1 U341 ( .A1(n398), .A2(n399), .ZN(n314) );
  NAND2_X1 U342 ( .A1(n400), .A2(n660), .ZN(n398) );
  NAND2_X1 U343 ( .A1(n515), .A2(n516), .ZN(n497) );
  NAND2_X1 U344 ( .A1(n81), .A2(n85), .ZN(n520) );
  INV_X1 U345 ( .A(n467), .ZN(n660) );
  INV_X1 U346 ( .A(n494), .ZN(n644) );
  INV_X1 U347 ( .A(n465), .ZN(n639) );
  NAND2_X1 U348 ( .A1(n98), .A2(n93), .ZN(n532) );
  AND2_X1 U349 ( .A1(n490), .A2(n489), .ZN(n481) );
  INV_X1 U350 ( .A(n113), .ZN(n592) );
  INV_X1 U351 ( .A(n484), .ZN(n643) );
  INV_X1 U352 ( .A(n102), .ZN(n590) );
  INV_X1 U353 ( .A(n375), .ZN(n579) );
  NOR2_X1 U354 ( .A1(B[61]), .A2(A[61]), .ZN(n71) );
  NOR2_X1 U355 ( .A1(n209), .A2(n208), .ZN(n207) );
  OR2_X1 U356 ( .A1(A[47]), .A2(B[47]), .ZN(n211) );
  NAND2_X1 U357 ( .A1(B[24]), .A2(A[24]), .ZN(n411) );
  NAND2_X1 U358 ( .A1(A[39]), .A2(B[39]), .ZN(n220) );
  NAND2_X1 U359 ( .A1(B[29]), .A2(A[29]), .ZN(n389) );
  NAND2_X1 U361 ( .A1(A[21]), .A2(B[21]), .ZN(n437) );
  NAND2_X1 U365 ( .A1(B[33]), .A2(A[33]), .ZN(n336) );
  NAND2_X1 U366 ( .A1(B[52]), .A2(A[52]), .ZN(n146) );
  NAND2_X1 U368 ( .A1(A[47]), .A2(B[47]), .ZN(n191) );
  NAND2_X1 U369 ( .A1(B[32]), .A2(A[32]), .ZN(n334) );
  NAND2_X1 U370 ( .A1(B[48]), .A2(A[48]), .ZN(n184) );
  OR2_X1 U371 ( .A1(B[28]), .A2(A[28]), .ZN(n380) );
  NAND2_X1 U372 ( .A1(B[20]), .A2(A[20]), .ZN(n438) );
  NAND2_X1 U373 ( .A1(B[36]), .A2(A[36]), .ZN(n307) );
  NAND2_X1 U374 ( .A1(B[62]), .A2(A[62]), .ZN(n107) );
  OR2_X1 U375 ( .A1(A[31]), .A2(B[31]), .ZN(n326) );
  OR2_X1 U377 ( .A1(B[24]), .A2(A[24]), .ZN(n413) );
  OR2_X1 U379 ( .A1(B[32]), .A2(A[32]), .ZN(n329) );
  NAND2_X1 U380 ( .A1(A[34]), .A2(B[34]), .ZN(n335) );
  NAND2_X1 U381 ( .A1(B[26]), .A2(A[26]), .ZN(n412) );
  NAND2_X1 U382 ( .A1(B[40]), .A2(A[40]), .ZN(n285) );
  NAND2_X1 U383 ( .A1(B[22]), .A2(A[22]), .ZN(n433) );
  NAND2_X1 U384 ( .A1(B[28]), .A2(A[28]), .ZN(n390) );
  OR2_X1 U385 ( .A1(B[27]), .A2(A[27]), .ZN(n360) );
  OR2_X1 U386 ( .A1(A[25]), .A2(B[25]), .ZN(n407) );
  NAND2_X1 U387 ( .A1(n171), .A2(n170), .ZN(n161) );
  AND2_X1 U388 ( .A1(n62), .A2(n63), .ZN(n283) );
  AND2_X1 U389 ( .A1(n303), .A2(n655), .ZN(n76) );
  OR2_X1 U390 ( .A1(B[62]), .A2(A[62]), .ZN(n113) );
  NAND2_X1 U391 ( .A1(B[27]), .A2(A[27]), .ZN(n421) );
  OR2_X1 U392 ( .A1(A[21]), .A2(B[21]), .ZN(n434) );
  NAND2_X1 U393 ( .A1(A[31]), .A2(B[31]), .ZN(n373) );
  OR2_X1 U394 ( .A1(A[23]), .A2(B[23]), .ZN(n431) );
  NAND2_X1 U395 ( .A1(B[63]), .A2(A[63]), .ZN(n106) );
  OR2_X1 U396 ( .A1(B[35]), .A2(A[35]), .ZN(n234) );
  OR2_X1 U397 ( .A1(A[47]), .A2(B[47]), .ZN(n30) );
  OR2_X1 U398 ( .A1(A[55]), .A2(B[55]), .ZN(n8) );
  OR2_X1 U399 ( .A1(B[63]), .A2(A[63]), .ZN(n102) );
  OR2_X1 U400 ( .A1(B[60]), .A2(A[60]), .ZN(n122) );
  OR2_X1 U401 ( .A1(B[18]), .A2(A[18]), .ZN(n457) );
  OR2_X1 U402 ( .A1(B[14]), .A2(A[14]), .ZN(n489) );
  OR2_X1 U403 ( .A1(B[19]), .A2(A[19]), .ZN(n458) );
  INV_X1 U404 ( .A(B[38]), .ZN(n655) );
  OR2_X1 U405 ( .A1(B[13]), .A2(A[13]), .ZN(n494) );
  OR2_X1 U406 ( .A1(B[17]), .A2(A[17]), .ZN(n465) );
  OR2_X1 U407 ( .A1(B[16]), .A2(A[16]), .ZN(n464) );
  OR2_X1 U408 ( .A1(B[15]), .A2(A[15]), .ZN(n490) );
  OR2_X1 U409 ( .A1(B[20]), .A2(A[20]), .ZN(n439) );
  INV_X1 U410 ( .A(B[41]), .ZN(n654) );
  OR2_X1 U411 ( .A1(B[6]), .A2(A[6]), .ZN(n93) );
  OR2_X1 U412 ( .A1(B[5]), .A2(A[5]), .ZN(n98) );
  OR2_X1 U413 ( .A1(B[10]), .A2(A[10]), .ZN(n521) );
  OR2_X1 U414 ( .A1(B[9]), .A2(A[9]), .ZN(n80) );
  OR2_X1 U415 ( .A1(B[11]), .A2(A[11]), .ZN(n515) );
  OR2_X1 U416 ( .A1(B[7]), .A2(A[7]), .ZN(n88) );
  OR2_X1 U417 ( .A1(B[8]), .A2(A[8]), .ZN(n84) );
  OR2_X1 U418 ( .A1(B[2]), .A2(A[2]), .ZN(n315) );
  OR2_X1 U419 ( .A1(B[12]), .A2(A[12]), .ZN(n493) );
  OR2_X1 U420 ( .A1(B[1]), .A2(A[1]), .ZN(n400) );
  OR2_X1 U421 ( .A1(B[4]), .A2(A[4]), .ZN(n130) );
  INV_X1 U422 ( .A(B[26]), .ZN(n657) );
  INV_X1 U423 ( .A(B[30]), .ZN(n656) );
  OR2_X1 U424 ( .A1(B[3]), .A2(A[3]), .ZN(n310) );
  OR2_X1 U425 ( .A1(B[0]), .A2(A[0]), .ZN(n534) );
  NAND2_X1 U426 ( .A1(B[1]), .A2(A[1]), .ZN(n399) );
  NAND2_X1 U427 ( .A1(B[8]), .A2(A[8]), .ZN(n85) );
  NAND2_X1 U428 ( .A1(B[12]), .A2(A[12]), .ZN(n486) );
  NAND2_X1 U429 ( .A1(B[14]), .A2(A[14]), .ZN(n488) );
  NAND2_X1 U430 ( .A1(B[13]), .A2(A[13]), .ZN(n487) );
  NAND2_X1 U431 ( .A1(B[17]), .A2(A[17]), .ZN(n462) );
  NAND2_X1 U432 ( .A1(B[6]), .A2(A[6]), .ZN(n90) );
  NAND2_X1 U433 ( .A1(B[16]), .A2(A[16]), .ZN(n461) );
  NAND2_X1 U434 ( .A1(B[18]), .A2(A[18]), .ZN(n463) );
  NAND2_X1 U435 ( .A1(B[9]), .A2(A[9]), .ZN(n81) );
  NAND2_X1 U436 ( .A1(B[2]), .A2(A[2]), .ZN(n312) );
  NAND2_X1 U437 ( .A1(B[0]), .A2(A[0]), .ZN(n467) );
  NAND2_X1 U438 ( .A1(B[4]), .A2(A[4]), .ZN(n129) );
  NAND2_X1 U439 ( .A1(B[5]), .A2(A[5]), .ZN(n97) );
  NAND2_X1 U440 ( .A1(B[10]), .A2(A[10]), .ZN(n518) );
  NAND2_X1 U441 ( .A1(B[19]), .A2(A[19]), .ZN(n456) );
  NAND2_X1 U442 ( .A1(B[3]), .A2(A[3]), .ZN(n311) );
  NAND2_X1 U443 ( .A1(B[7]), .A2(A[7]), .ZN(n89) );
  NAND2_X1 U444 ( .A1(B[15]), .A2(A[15]), .ZN(n484) );
  NAND2_X1 U445 ( .A1(B[11]), .A2(A[11]), .ZN(n519) );
  NAND2_X1 U446 ( .A1(A[38]), .A2(B[38]), .ZN(n318) );
  OR2_X1 U447 ( .A1(B[38]), .A2(A[38]), .ZN(n63) );
  NOR3_X1 U448 ( .A1(n630), .A2(n348), .A3(n19), .ZN(n224) );
  AOI21_X1 U449 ( .B1(n334), .B2(n233), .A(n342), .ZN(n339) );
  OAI21_X1 U450 ( .B1(n572), .B2(n71), .A(n110), .ZN(n115) );
  AOI22_X1 U451 ( .A1(A[31]), .A2(B[31]), .B1(n371), .B2(n582), .ZN(n354) );
  AOI21_X1 U452 ( .B1(n656), .B2(n581), .A(n579), .ZN(n371) );
  NAND2_X1 U453 ( .A1(B[54]), .A2(A[54]), .ZN(n148) );
  XNOR2_X1 U454 ( .A(n343), .B(n344), .ZN(SUM[34]) );
  XNOR2_X1 U455 ( .A(n2), .B(n387), .ZN(SUM[31]) );
  OAI21_X1 U456 ( .B1(n11), .B2(n388), .A(n386), .ZN(n387) );
  NAND2_X1 U457 ( .A1(A[43]), .A2(B[43]), .ZN(n257) );
  AND2_X1 U458 ( .A1(B[43]), .A2(n542), .ZN(n77) );
  OR2_X1 U459 ( .A1(B[43]), .A2(A[43]), .ZN(n212) );
  NAND2_X1 U460 ( .A1(B[49]), .A2(A[49]), .ZN(n163) );
  AND2_X1 U461 ( .A1(B[49]), .A2(A[49]), .ZN(n72) );
  NAND2_X1 U462 ( .A1(B[61]), .A2(A[61]), .ZN(n110) );
  OAI21_X1 U463 ( .B1(n51), .B2(n576), .A(n410), .ZN(n420) );
  OAI21_X1 U464 ( .B1(n51), .B2(n576), .A(n410), .ZN(n31) );
  INV_X1 U465 ( .A(n234), .ZN(n630) );
  NAND2_X1 U466 ( .A1(n56), .A2(n234), .ZN(n325) );
  NAND2_X1 U467 ( .A1(B[35]), .A2(n543), .ZN(n222) );
  OR2_X1 U468 ( .A1(A[35]), .A2(B[35]), .ZN(n337) );
  NAND4_X1 U469 ( .A1(n354), .A2(n353), .A3(n352), .A4(n355), .ZN(n324) );
  NAND4_X1 U470 ( .A1(n354), .A2(n353), .A3(n352), .A4(n355), .ZN(n29) );
  NAND2_X1 U471 ( .A1(n181), .A2(n180), .ZN(n179) );
  NAND2_X1 U472 ( .A1(B[44]), .A2(A[44]), .ZN(n201) );
  NAND2_X1 U473 ( .A1(n420), .A2(n409), .ZN(n419) );
  AND2_X1 U474 ( .A1(n139), .A2(n140), .ZN(n141) );
  AOI21_X1 U475 ( .B1(n273), .B2(n272), .A(n274), .ZN(n271) );
  NAND2_X1 U476 ( .A1(net489128), .A2(n594), .ZN(net489130) );
  INV_X1 U477 ( .A(net537531), .ZN(n594) );
  NAND2_X1 U478 ( .A1(B[58]), .A2(A[58]), .ZN(net489105) );
  INV_X1 U479 ( .A(n122), .ZN(n588) );
  NAND2_X1 U480 ( .A1(n161), .A2(n169), .ZN(n136) );
  NAND2_X1 U481 ( .A1(A[51]), .A2(B[51]), .ZN(n160) );
  OR2_X1 U482 ( .A1(A[51]), .A2(B[51]), .ZN(n172) );
  OR2_X1 U483 ( .A1(A[51]), .A2(B[51]), .ZN(n59) );
  AOI21_X1 U484 ( .B1(n141), .B2(n142), .A(n599), .ZN(n132) );
  INV_X1 U485 ( .A(n144), .ZN(n599) );
  INV_X1 U486 ( .A(A[38]), .ZN(n621) );
  NAND2_X1 U487 ( .A1(n147), .A2(n138), .ZN(n165) );
  AND2_X1 U488 ( .A1(n137), .A2(n138), .ZN(n135) );
  NAND2_X1 U489 ( .A1(n304), .A2(n76), .ZN(n62) );
  OAI211_X1 U490 ( .C1(B[30]), .C2(A[30]), .A(n380), .B(n375), .ZN(n25) );
  NAND2_X1 U491 ( .A1(A[30]), .A2(B[30]), .ZN(n386) );
  INV_X1 U492 ( .A(A[30]), .ZN(n581) );
  AND2_X1 U493 ( .A1(A[57]), .A2(B[57]), .ZN(net537531) );
  NAND2_X1 U494 ( .A1(A[46]), .A2(B[46]), .ZN(n202) );
  NAND2_X1 U495 ( .A1(n111), .A2(n122), .ZN(n124) );
  OAI21_X1 U496 ( .B1(n573), .B2(n588), .A(n111), .ZN(n121) );
  OAI211_X1 U497 ( .C1(n573), .C2(n588), .A(n110), .B(n111), .ZN(n104) );
  XNOR2_X1 U498 ( .A(n114), .B(n10), .ZN(SUM[63]) );
  AND2_X1 U499 ( .A1(n106), .A2(n102), .ZN(n10) );
  INV_X1 U500 ( .A(n258), .ZN(n601) );
  AND2_X1 U501 ( .A1(n258), .A2(n7), .ZN(n64) );
  AND2_X1 U502 ( .A1(n257), .A2(n258), .ZN(n256) );
  AND2_X1 U503 ( .A1(B[59]), .A2(A[59]), .ZN(n73) );
  XNOR2_X1 U504 ( .A(n115), .B(n117), .ZN(SUM[62]) );
  NAND2_X1 U505 ( .A1(n113), .A2(n107), .ZN(n117) );
  XNOR2_X1 U506 ( .A(n52), .B(n321), .ZN(SUM[37]) );
  NAND4_X1 U507 ( .A1(n193), .A2(n36), .A3(n190), .A4(n191), .ZN(n170) );
  NAND4_X1 U508 ( .A1(n193), .A2(n190), .A3(n192), .A4(n191), .ZN(n189) );
  XNOR2_X1 U509 ( .A(net489114), .B(n131), .ZN(SUM[59]) );
  OAI21_X1 U510 ( .B1(n575), .B2(n277), .A(n278), .ZN(n273) );
  XNOR2_X1 U511 ( .A(n124), .B(n123), .ZN(SUM[60]) );
  NOR2_X1 U512 ( .A1(n589), .A2(n71), .ZN(n119) );
  AND2_X1 U513 ( .A1(n162), .A2(n559), .ZN(n54) );
  AND2_X1 U514 ( .A1(n164), .A2(n559), .ZN(n5) );
  NAND2_X1 U515 ( .A1(n164), .A2(n173), .ZN(n185) );
  OR2_X1 U516 ( .A1(n205), .A2(n9), .ZN(n53) );
  NAND2_X1 U517 ( .A1(n9), .A2(n249), .ZN(n248) );
  NAND2_X1 U518 ( .A1(B[41]), .A2(A[41]), .ZN(n286) );
  INV_X1 U519 ( .A(A[41]), .ZN(n616) );
  OAI211_X1 U520 ( .C1(n555), .C2(n334), .A(n335), .B(n336), .ZN(n332) );
  NAND2_X1 U521 ( .A1(net489125), .A2(net489103), .ZN(net489131) );
  NAND2_X1 U522 ( .A1(net489099), .A2(net489103), .ZN(net489134) );
  NAND4_X1 U523 ( .A1(n439), .A2(n434), .A3(n435), .A4(n431), .ZN(n368) );
  NAND2_X1 U524 ( .A1(n434), .A2(n437), .ZN(n448) );
  AND3_X1 U525 ( .A1(n436), .A2(n435), .A3(n434), .ZN(n429) );
  INV_X1 U526 ( .A(n434), .ZN(n633) );
  NAND4_X1 U529 ( .A1(n228), .A2(n566), .A3(n230), .A4(n554), .ZN(n223) );
  NAND2_X1 U530 ( .A1(n303), .A2(n229), .ZN(n321) );
  INV_X1 U531 ( .A(n229), .ZN(n620) );
  NAND2_X1 U532 ( .A1(n229), .A2(n604), .ZN(n304) );
  NAND2_X1 U536 ( .A1(B[55]), .A2(A[55]), .ZN(n144) );
  OR2_X1 U537 ( .A1(A[55]), .A2(B[55]), .ZN(n139) );
  INV_X1 U539 ( .A(n18), .ZN(n584) );
  NAND2_X1 U540 ( .A1(B[60]), .A2(A[60]), .ZN(n111) );
  NAND2_X1 U541 ( .A1(n132), .A2(n133), .ZN(net489093) );
  XNOR2_X1 U542 ( .A(n295), .B(n296), .ZN(SUM[41]) );
  NAND2_X1 U543 ( .A1(n211), .A2(n210), .ZN(n209) );
  NAND2_X1 U544 ( .A1(n188), .A2(n184), .ZN(n187) );
  AOI21_X1 U545 ( .B1(net489120), .B2(net489106), .A(n596), .ZN(net489114) );
  XNOR2_X1 U546 ( .A(net489122), .B(net489120), .ZN(SUM[58]) );
  AOI21_X1 U547 ( .B1(n288), .B2(n289), .A(n617), .ZN(n287) );
  NAND2_X1 U548 ( .A1(n432), .A2(n431), .ZN(n440) );
  NAND2_X1 U549 ( .A1(n432), .A2(n433), .ZN(n430) );
  NOR2_X1 U551 ( .A1(n561), .A2(n614), .ZN(n249) );
  AOI21_X1 U552 ( .B1(n18), .B2(n175), .A(n585), .ZN(n169) );
  AND2_X1 U554 ( .A1(n59), .A2(n559), .ZN(n18) );
  INV_X1 U555 ( .A(n160), .ZN(n585) );
  XNOR2_X1 U558 ( .A(n166), .B(n165), .ZN(SUM[53]) );
  XNOR2_X1 U559 ( .A(n319), .B(n320), .ZN(SUM[38]) );
  AOI21_X1 U560 ( .B1(n319), .B2(n230), .A(n622), .ZN(n22) );
  OAI21_X1 U561 ( .B1(n20), .B2(n620), .A(n303), .ZN(n319) );
  INV_X1 U562 ( .A(n549), .ZN(n574) );
  AOI21_X1 U563 ( .B1(n28), .B2(n228), .A(n604), .ZN(n20) );
  XNOR2_X1 U564 ( .A(n150), .B(n151), .ZN(SUM[55]) );
  INV_X1 U565 ( .A(n121), .ZN(n572) );
  NAND2_X1 U567 ( .A1(n125), .A2(net489091), .ZN(n123) );
  AOI21_X1 U568 ( .B1(n126), .B2(net489101), .A(n73), .ZN(n125) );
  NOR2_X1 U569 ( .A1(n73), .A2(n74), .ZN(n131) );
  NOR2_X1 U570 ( .A1(n595), .A2(n74), .ZN(n126) );
  XNOR2_X1 U571 ( .A(n235), .B(n65), .ZN(SUM[47]) );
  XNOR2_X1 U572 ( .A(n186), .B(n54), .ZN(SUM[50]) );
  AOI21_X1 U573 ( .B1(n187), .B2(n164), .A(n72), .ZN(n186) );
  NOR2_X1 U576 ( .A1(n271), .A2(n601), .ZN(n268) );
  NAND2_X1 U577 ( .A1(A[37]), .A2(B[37]), .ZN(n303) );
  XNOR2_X1 U578 ( .A(net489130), .B(net489131), .ZN(SUM[57]) );
  AOI21_X1 U579 ( .B1(n382), .B2(n403), .A(n12), .ZN(n404) );
  INV_X1 U581 ( .A(n367), .ZN(n631) );
  XNOR2_X1 U582 ( .A(n427), .B(n403), .ZN(SUM[24]) );
  NAND2_X1 U583 ( .A1(n403), .A2(n413), .ZN(n426) );
  AOI21_X1 U585 ( .B1(n403), .B2(n413), .A(n577), .ZN(n51) );
  NAND2_X1 U586 ( .A1(A[23]), .A2(B[23]), .ZN(n432) );
  XNOR2_X1 U587 ( .A(n156), .B(n157), .ZN(SUM[54]) );
  NAND2_X1 U589 ( .A1(B[53]), .A2(A[53]), .ZN(n147) );
  XNOR2_X1 U590 ( .A(n338), .B(n50), .ZN(SUM[35]) );
  NAND2_X1 U591 ( .A1(n29), .A2(n548), .ZN(n233) );
  NAND2_X1 U592 ( .A1(n548), .A2(n29), .ZN(n19) );
  AOI21_X1 U593 ( .B1(net489128), .B2(n597), .A(net537531), .ZN(net489126) );
  INV_X1 U597 ( .A(net489103), .ZN(n597) );
  OAI21_X1 U598 ( .B1(n593), .B2(net489125), .A(net489126), .ZN(net489120) );
  NAND2_X1 U600 ( .A1(net489093), .A2(net489099), .ZN(net489125) );
  AOI21_X1 U601 ( .B1(n135), .B2(n154), .A(n155), .ZN(n156) );
  NAND2_X1 U602 ( .A1(n155), .A2(n140), .ZN(n152) );
  XNOR2_X1 U603 ( .A(n287), .B(n64), .ZN(SUM[42]) );
  NAND2_X1 U604 ( .A1(A[50]), .A2(B[50]), .ZN(n162) );
  XNOR2_X1 U605 ( .A(n252), .B(n297), .ZN(SUM[40]) );
  NAND2_X1 U606 ( .A1(n226), .A2(n252), .ZN(n42) );
  AOI21_X1 U607 ( .B1(n252), .B2(n265), .A(n618), .ZN(n295) );
  NAND2_X1 U608 ( .A1(B[56]), .A2(A[56]), .ZN(net489103) );
  XNOR2_X1 U609 ( .A(n556), .B(net489134), .ZN(SUM[56]) );
  NAND2_X1 U610 ( .A1(A[42]), .A2(B[42]), .ZN(n258) );
  OR2_X1 U611 ( .A1(A[42]), .A2(B[42]), .ZN(n259) );
  XNOR2_X1 U612 ( .A(n242), .B(n243), .ZN(SUM[46]) );
  XNOR2_X1 U613 ( .A(n572), .B(n119), .ZN(SUM[61]) );
  NAND4_X1 U614 ( .A1(B[27]), .A2(n414), .A3(n413), .A4(n407), .ZN(n362) );
  NAND4_X1 U615 ( .A1(n414), .A2(n407), .A3(A[27]), .A4(n413), .ZN(n363) );
  NAND2_X1 U616 ( .A1(n407), .A2(n410), .ZN(n425) );
  INV_X1 U617 ( .A(n407), .ZN(n576) );
  NAND2_X1 U618 ( .A1(B[25]), .A2(A[25]), .ZN(n410) );
  OAI211_X1 U619 ( .C1(n593), .C2(net489103), .A(n594), .B(net489105), .ZN(
        net489101) );
  NAND2_X1 U620 ( .A1(net489106), .A2(net489105), .ZN(net489122) );
  INV_X1 U621 ( .A(net489105), .ZN(n596) );
  INV_X1 U622 ( .A(n110), .ZN(n589) );
  NOR2_X1 U623 ( .A1(B[59]), .A2(A[59]), .ZN(n74) );
endmodule


module RCA_NBIT64_6 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_6_DW01_add_8 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_5_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net487998, net487988, net487987, net487986, net487985, net487981,
         net487964, net487952, net487950, net487948, net487943, net487940,
         net487918, net487915, net487913, net487908, net487907, net538236,
         net487929, net487910, net487930, net487920, net487984, net487983,
         net487939, net487938, net487933, net487931, net487921, net487919, n3,
         n5, n7, n9, n10, n13, n14, n15, n16, n17, n18, n19, n24, n25, n26,
         n27, n34, n36, n37, n39, n46, n47, n52, n53, n54, n55, n56, n59, n60,
         n61, n62, n63, n64, n65, n67, n68, n69, n70, n71, n72, n74, n75, n76,
         n78, n79, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n116, n117, n120, n121, n122, n123,
         n124, n125, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n157, n158, n159, n160,
         n161, n162, n163, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n179, n180, n181, n182, n184, n185,
         n186, n188, n189, n190, n191, n193, n197, n198, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n219, n220, n221, n222, n223, n224, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n238, n241, n242, n243,
         n244, n245, n246, n249, n250, n251, n252, n253, n254, n256, n257,
         n258, n259, n260, n262, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n274, n275, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n293, n295, n298,
         n299, n300, n303, n304, n305, n308, n309, n310, n311, n312, n313,
         n314, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n346, n347, n348, n349, n350, n352, n353,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n368,
         n370, n371, n372, n373, n374, n375, n377, n378, n379, n380, n381,
         n382, n383, n385, n386, n387, n388, n389, n390, n392, n393, n394,
         n395, n397, n399, n402, n403, n404, n406, n407, n408, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n421, n422, n423, n424,
         n425, n426, n428, n430, n431, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n451, n452, n453, n454, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n473, n474, n476,
         n477, n481, n482, n483, n484, n485, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n502, n503,
         n504, n505, n506, n507, n508, n510, n512, n513, n514, n515, n516,
         n519, n520, n521, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n555,
         n556, n557, n558, n560, n562, n563, n564, n565, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686;

  OR2_X2 U25 ( .A1(A[54]), .A2(B[54]), .ZN(net487981) );
  NAND3_X1 U50 ( .A1(n350), .A2(n46), .A3(n574), .ZN(n27) );
  NAND3_X1 U59 ( .A1(n65), .A2(n575), .A3(n270), .ZN(n304) );
  NAND3_X1 U62 ( .A1(n327), .A2(n328), .A3(n323), .ZN(n317) );
  NAND3_X1 U68 ( .A1(n70), .A2(n54), .A3(n175), .ZN(n59) );
  OR2_X2 U85 ( .A1(A[56]), .A2(B[56]), .ZN(net487913) );
  OR2_X2 U119 ( .A1(A[39]), .A2(B[39]), .ZN(n270) );
  NAND3_X1 U129 ( .A1(n143), .A2(n144), .A3(n145), .ZN(n56) );
  OR2_X2 U145 ( .A1(B[48]), .A2(A[48]), .ZN(n198) );
  NAND3_X1 U148 ( .A1(n433), .A2(n581), .A3(n15), .ZN(n394) );
  NAND3_X1 U151 ( .A1(n61), .A2(n169), .A3(n14), .ZN(n206) );
  OR2_X2 U156 ( .A1(A[44]), .A2(B[44]), .ZN(n244) );
  OR2_X2 U158 ( .A1(A[34]), .A2(B[34]), .ZN(n237) );
  OR2_X2 U370 ( .A1(A[37]), .A2(B[37]), .ZN(n268) );
  OR2_X2 U379 ( .A1(B[36]), .A2(A[36]), .ZN(n267) );
  OR2_X2 U390 ( .A1(B[40]), .A2(A[40]), .ZN(n291) );
  NAND3_X1 U563 ( .A1(n158), .A2(net487981), .A3(n25), .ZN(n147) );
  NAND3_X1 U566 ( .A1(n167), .A2(n168), .A3(n205), .ZN(n166) );
  NAND3_X1 U573 ( .A1(n157), .A2(n54), .A3(n181), .ZN(n193) );
  NAND3_X1 U577 ( .A1(n154), .A2(n181), .A3(n54), .ZN(n197) );
  NAND3_X1 U578 ( .A1(A[48]), .A2(B[48]), .A3(n185), .ZN(n167) );
  NAND3_X1 U579 ( .A1(n204), .A2(n206), .A3(n205), .ZN(n203) );
  NAND3_X1 U580 ( .A1(n169), .A2(n208), .A3(n207), .ZN(n204) );
  NAND3_X1 U581 ( .A1(n168), .A2(n212), .A3(n213), .ZN(n211) );
  NAND3_X1 U582 ( .A1(n61), .A2(n207), .A3(n198), .ZN(n213) );
  NAND3_X1 U587 ( .A1(n630), .A2(n574), .A3(n238), .ZN(n234) );
  NAND3_X1 U589 ( .A1(n262), .A2(n69), .A3(n253), .ZN(n260) );
  NAND3_X1 U594 ( .A1(n290), .A2(n289), .A3(n288), .ZN(n286) );
  NAND3_X1 U601 ( .A1(n252), .A2(n69), .A3(n300), .ZN(n299) );
  NAND3_X1 U607 ( .A1(n258), .A2(n257), .A3(n304), .ZN(n311) );
  NAND3_X1 U609 ( .A1(n268), .A2(n324), .A3(n269), .ZN(n323) );
  NAND3_X1 U618 ( .A1(n237), .A2(n352), .A3(n353), .ZN(n364) );
  NAND3_X1 U623 ( .A1(n390), .A2(n389), .A3(n388), .ZN(n379) );
  NAND3_X1 U640 ( .A1(n435), .A2(n436), .A3(n437), .ZN(n434) );
  NAND3_X1 U641 ( .A1(n438), .A2(n439), .A3(n440), .ZN(n435) );
  NAND3_X1 U666 ( .A1(n543), .A2(n544), .A3(n545), .ZN(n542) );
  NAND3_X1 U667 ( .A1(n546), .A2(n86), .A3(n547), .ZN(n543) );
  CLKBUF_X1 U2 ( .A(A[54]), .Z(n568) );
  AND2_X1 U3 ( .A1(n571), .A2(B[51]), .ZN(n569) );
  OR2_X1 U4 ( .A1(B[55]), .A2(A[55]), .ZN(net487964) );
  OR2_X1 U5 ( .A1(B[52]), .A2(A[52]), .ZN(n25) );
  AND2_X1 U6 ( .A1(net487984), .A2(net487983), .ZN(net538236) );
  AND2_X1 U7 ( .A1(n560), .A2(n493), .ZN(SUM[0]) );
  OR2_X1 U8 ( .A1(B[59]), .A2(A[59]), .ZN(net487910) );
  CLKBUF_X1 U9 ( .A(A[53]), .Z(n570) );
  CLKBUF_X1 U10 ( .A(A[51]), .Z(n571) );
  AND2_X1 U11 ( .A1(net487918), .A2(net487938), .ZN(n572) );
  INV_X1 U12 ( .A(B[45]), .ZN(n585) );
  XNOR2_X1 U13 ( .A(n573), .B(n36), .ZN(SUM[39]) );
  AND2_X1 U14 ( .A1(n270), .A2(n327), .ZN(n573) );
  OR2_X1 U15 ( .A1(A[38]), .A2(B[38]), .ZN(n576) );
  OR2_X1 U16 ( .A1(A[43]), .A2(B[43]), .ZN(n253) );
  NAND3_X1 U17 ( .A1(net487919), .A2(net487939), .A3(n572), .ZN(net487933) );
  CLKBUF_X1 U18 ( .A(n237), .Z(n574) );
  NAND2_X1 U19 ( .A1(n26), .A2(n27), .ZN(n575) );
  NOR2_X1 U20 ( .A1(A[42]), .A2(B[42]), .ZN(n293) );
  AND3_X1 U21 ( .A1(n327), .A2(n328), .A3(n323), .ZN(n577) );
  OR2_X1 U22 ( .A1(A[38]), .A2(B[38]), .ZN(n269) );
  OR2_X1 U23 ( .A1(B[57]), .A2(A[57]), .ZN(n578) );
  OR2_X1 U24 ( .A1(B[57]), .A2(A[57]), .ZN(net487921) );
  NAND2_X1 U26 ( .A1(n65), .A2(n9), .ZN(n579) );
  INV_X1 U27 ( .A(n591), .ZN(n580) );
  OR2_X1 U28 ( .A1(B[26]), .A2(A[26]), .ZN(n581) );
  OR2_X1 U29 ( .A1(A[26]), .A2(B[26]), .ZN(n440) );
  OR2_X1 U30 ( .A1(A[49]), .A2(B[49]), .ZN(n207) );
  OAI21_X1 U31 ( .B1(n601), .B2(n654), .A(n386), .ZN(n582) );
  OR2_X1 U32 ( .A1(B[50]), .A2(A[50]), .ZN(n54) );
  AND2_X1 U33 ( .A1(n298), .A2(n299), .ZN(n583) );
  AND2_X1 U34 ( .A1(n576), .A2(n330), .ZN(n65) );
  OR2_X1 U35 ( .A1(B[41]), .A2(A[41]), .ZN(n254) );
  OR2_X1 U36 ( .A1(B[41]), .A2(A[41]), .ZN(n69) );
  OR2_X1 U37 ( .A1(n585), .A2(n644), .ZN(n227) );
  AND2_X1 U38 ( .A1(n244), .A2(n245), .ZN(n584) );
  AND3_X1 U39 ( .A1(n246), .A2(n16), .A3(n584), .ZN(n243) );
  AND2_X1 U40 ( .A1(n644), .A2(n585), .ZN(n228) );
  AND2_X1 U41 ( .A1(n55), .A2(n167), .ZN(n586) );
  NAND2_X1 U42 ( .A1(n587), .A2(n174), .ZN(n588) );
  AND2_X1 U43 ( .A1(n157), .A2(net487981), .ZN(n587) );
  NOR2_X1 U44 ( .A1(n588), .A2(n589), .ZN(n159) );
  AND2_X1 U45 ( .A1(n59), .A2(n163), .ZN(n589) );
  AND2_X2 U46 ( .A1(n624), .A2(n681), .ZN(n71) );
  NAND2_X1 U47 ( .A1(n158), .A2(n157), .ZN(n590) );
  NOR2_X1 U48 ( .A1(B[58]), .A2(A[58]), .ZN(n591) );
  OR2_X1 U49 ( .A1(A[45]), .A2(B[45]), .ZN(n245) );
  AND2_X1 U51 ( .A1(n644), .A2(n585), .ZN(n592) );
  NOR2_X1 U52 ( .A1(n592), .A2(n282), .ZN(n280) );
  XNOR2_X1 U53 ( .A(n593), .B(n594), .ZN(SUM[52]) );
  NAND3_X1 U54 ( .A1(n197), .A2(n180), .A3(n59), .ZN(n593) );
  NAND2_X1 U55 ( .A1(net487986), .A2(n25), .ZN(n594) );
  OR2_X1 U56 ( .A1(B[43]), .A2(A[43]), .ZN(n305) );
  INV_X1 U57 ( .A(n444), .ZN(n657) );
  INV_X1 U58 ( .A(n476), .ZN(n662) );
  AOI21_X1 U60 ( .B1(n142), .B2(net487940), .A(net487950), .ZN(net487948) );
  NOR2_X1 U61 ( .A1(n622), .A2(n623), .ZN(n79) );
  OAI21_X1 U63 ( .B1(n662), .B2(n413), .A(n399), .ZN(n444) );
  AOI21_X1 U64 ( .B1(n658), .B2(n397), .A(n656), .ZN(n393) );
  INV_X1 U65 ( .A(n399), .ZN(n656) );
  OAI21_X1 U66 ( .B1(n5), .B2(n342), .A(n343), .ZN(n24) );
  NAND2_X1 U67 ( .A1(n150), .A2(n146), .ZN(net487940) );
  NOR2_X1 U69 ( .A1(n623), .A2(n147), .ZN(n150) );
  NAND2_X1 U70 ( .A1(n579), .A2(n258), .ZN(n289) );
  INV_X1 U71 ( .A(n235), .ZN(n633) );
  INV_X1 U72 ( .A(n313), .ZN(n639) );
  INV_X1 U73 ( .A(n188), .ZN(n608) );
  AND2_X1 U74 ( .A1(n74), .A2(n577), .ZN(n319) );
  INV_X1 U75 ( .A(n373), .ZN(n630) );
  OAI21_X1 U76 ( .B1(n684), .B2(n528), .A(n525), .ZN(n89) );
  OAI21_X1 U77 ( .B1(n668), .B2(n411), .A(n663), .ZN(n476) );
  INV_X1 U78 ( .A(n397), .ZN(n663) );
  INV_X1 U79 ( .A(n402), .ZN(n668) );
  AOI21_X1 U80 ( .B1(n524), .B2(n525), .A(n526), .ZN(n521) );
  NAND2_X1 U81 ( .A1(n676), .A2(n527), .ZN(n524) );
  INV_X1 U82 ( .A(n528), .ZN(n676) );
  NAND2_X1 U83 ( .A1(n540), .A2(n523), .ZN(n538) );
  NAND2_X1 U84 ( .A1(n672), .A2(n89), .ZN(n540) );
  INV_X1 U86 ( .A(n526), .ZN(n672) );
  INV_X1 U87 ( .A(n394), .ZN(n603) );
  INV_X1 U88 ( .A(n413), .ZN(n658) );
  INV_X1 U89 ( .A(n527), .ZN(n684) );
  INV_X1 U90 ( .A(n411), .ZN(n664) );
  NOR2_X1 U91 ( .A1(n106), .A2(n620), .ZN(SUM[64]) );
  INV_X1 U92 ( .A(n406), .ZN(n652) );
  INV_X1 U93 ( .A(n523), .ZN(n673) );
  NAND2_X1 U94 ( .A1(n69), .A2(n256), .ZN(n321) );
  NAND2_X1 U95 ( .A1(n270), .A2(n291), .ZN(n320) );
  NOR2_X1 U96 ( .A1(n647), .A2(n82), .ZN(n275) );
  INV_X1 U97 ( .A(n229), .ZN(n647) );
  INV_X1 U98 ( .A(n223), .ZN(n646) );
  AND2_X1 U99 ( .A1(n438), .A2(n443), .ZN(n15) );
  XOR2_X1 U100 ( .A(n56), .B(n595), .Z(SUM[57]) );
  AND2_X1 U101 ( .A1(n578), .A2(net487919), .ZN(n595) );
  NOR2_X1 U102 ( .A1(n642), .A2(n641), .ZN(n60) );
  AOI22_X1 U103 ( .A1(n281), .A2(n253), .B1(n635), .B2(n289), .ZN(n295) );
  INV_X1 U104 ( .A(n287), .ZN(n641) );
  NOR2_X1 U105 ( .A1(n645), .A2(n83), .ZN(n284) );
  NOR2_X1 U106 ( .A1(n583), .A2(n282), .ZN(n285) );
  AOI211_X1 U107 ( .C1(n258), .C2(n259), .A(n260), .B(n643), .ZN(n241) );
  INV_X1 U108 ( .A(n291), .ZN(n643) );
  NAND2_X1 U109 ( .A1(n633), .A2(n264), .ZN(n259) );
  NAND2_X1 U110 ( .A1(n421), .A2(n386), .ZN(n428) );
  NAND2_X1 U111 ( .A1(n209), .A2(n198), .ZN(n219) );
  NAND2_X1 U112 ( .A1(n267), .A2(n326), .ZN(n349) );
  NAND2_X1 U113 ( .A1(n581), .A2(n436), .ZN(n449) );
  AND2_X1 U114 ( .A1(n251), .A2(n253), .ZN(n309) );
  AOI21_X1 U115 ( .B1(n310), .B2(n311), .A(n312), .ZN(n308) );
  NOR2_X1 U116 ( .A1(n293), .A2(n313), .ZN(n310) );
  NOR2_X1 U117 ( .A1(n627), .A2(n626), .ZN(n216) );
  INV_X1 U118 ( .A(n207), .ZN(n626) );
  XNOR2_X1 U120 ( .A(n452), .B(n451), .ZN(SUM[25]) );
  NAND2_X1 U121 ( .A1(n438), .A2(n441), .ZN(n452) );
  NAND2_X1 U122 ( .A1(n453), .A2(n442), .ZN(n451) );
  NAND2_X1 U123 ( .A1(n39), .A2(net487910), .ZN(net487929) );
  NAND2_X1 U124 ( .A1(n606), .A2(n207), .ZN(n212) );
  XNOR2_X1 U125 ( .A(n314), .B(n63), .ZN(SUM[42]) );
  NOR2_X1 U126 ( .A1(n293), .A2(n637), .ZN(n63) );
  AOI21_X1 U127 ( .B1(n639), .B2(n311), .A(n640), .ZN(n314) );
  INV_X1 U128 ( .A(n256), .ZN(n640) );
  AOI21_X1 U130 ( .B1(n24), .B2(n576), .A(n634), .ZN(n36) );
  INV_X1 U131 ( .A(n328), .ZN(n634) );
  XNOR2_X1 U132 ( .A(n363), .B(n362), .ZN(SUM[35]) );
  NAND2_X1 U133 ( .A1(n266), .A2(n361), .ZN(n362) );
  OAI21_X1 U134 ( .B1(n364), .B2(n372), .A(n365), .ZN(n363) );
  OAI21_X1 U135 ( .B1(n17), .B2(n456), .A(n457), .ZN(n399) );
  AND3_X1 U136 ( .A1(n460), .A2(n461), .A3(n462), .ZN(n17) );
  NAND2_X1 U137 ( .A1(n463), .A2(n464), .ZN(n461) );
  NAND4_X1 U138 ( .A1(n378), .A2(n379), .A3(n380), .A4(n381), .ZN(n46) );
  XNOR2_X1 U139 ( .A(n377), .B(n46), .ZN(SUM[32]) );
  NAND2_X1 U140 ( .A1(n352), .A2(n359), .ZN(n377) );
  XNOR2_X1 U141 ( .A(n431), .B(n47), .ZN(SUM[28]) );
  NAND2_X1 U142 ( .A1(n412), .A2(n385), .ZN(n431) );
  OAI21_X1 U143 ( .B1(n657), .B2(n394), .A(n395), .ZN(n47) );
  XNOR2_X1 U144 ( .A(n454), .B(n444), .ZN(SUM[24]) );
  NAND2_X1 U146 ( .A1(n443), .A2(n442), .ZN(n454) );
  XNOR2_X1 U147 ( .A(n374), .B(n375), .ZN(SUM[33]) );
  AOI21_X1 U149 ( .B1(n352), .B2(n230), .A(n629), .ZN(n374) );
  NOR2_X1 U150 ( .A1(n650), .A2(n651), .ZN(n375) );
  INV_X1 U152 ( .A(n353), .ZN(n651) );
  XNOR2_X1 U153 ( .A(n474), .B(n473), .ZN(SUM[21]) );
  NAND2_X1 U154 ( .A1(n460), .A2(n463), .ZN(n474) );
  NAND2_X1 U155 ( .A1(n237), .A2(n368), .ZN(n370) );
  XNOR2_X1 U157 ( .A(n75), .B(n322), .ZN(SUM[40]) );
  NAND2_X1 U159 ( .A1(n291), .A2(n257), .ZN(n322) );
  NAND2_X1 U160 ( .A1(n304), .A2(n258), .ZN(n75) );
  XNOR2_X1 U161 ( .A(n341), .B(n67), .ZN(SUM[38]) );
  NAND2_X1 U162 ( .A1(n328), .A2(n576), .ZN(n67) );
  OAI21_X1 U163 ( .B1(n5), .B2(n342), .A(n343), .ZN(n341) );
  XNOR2_X1 U164 ( .A(n415), .B(n414), .ZN(SUM[31]) );
  NAND2_X1 U165 ( .A1(n381), .A2(n392), .ZN(n414) );
  NAND2_X1 U166 ( .A1(n608), .A2(n54), .ZN(n186) );
  AOI21_X1 U167 ( .B1(n650), .B2(n237), .A(n631), .ZN(n365) );
  INV_X1 U168 ( .A(n368), .ZN(n631) );
  OAI21_X1 U169 ( .B1(n602), .B2(n604), .A(n385), .ZN(n422) );
  INV_X1 U170 ( .A(n412), .ZN(n604) );
  INV_X1 U171 ( .A(n430), .ZN(n602) );
  OAI21_X1 U172 ( .B1(n394), .B2(n657), .A(n395), .ZN(n430) );
  OAI21_X1 U173 ( .B1(n19), .B2(n655), .A(n441), .ZN(n448) );
  INV_X1 U174 ( .A(n438), .ZN(n655) );
  AND2_X1 U175 ( .A1(n453), .A2(n442), .ZN(n19) );
  XNOR2_X1 U176 ( .A(n121), .B(n122), .ZN(SUM[63]) );
  NAND2_X1 U177 ( .A1(n113), .A2(n123), .ZN(n121) );
  NAND2_X1 U178 ( .A1(n112), .A2(n108), .ZN(n122) );
  XNOR2_X1 U179 ( .A(n347), .B(n346), .ZN(SUM[37]) );
  NAND2_X1 U180 ( .A1(n348), .A2(n326), .ZN(n347) );
  OAI21_X1 U181 ( .B1(n293), .B2(n256), .A(n303), .ZN(n312) );
  OAI21_X1 U182 ( .B1(n249), .B2(n250), .A(n251), .ZN(n242) );
  AOI21_X1 U183 ( .B1(n300), .B2(n69), .A(n637), .ZN(n249) );
  NAND2_X1 U184 ( .A1(n252), .A2(n253), .ZN(n250) );
  NAND2_X1 U185 ( .A1(n298), .A2(n299), .ZN(n281) );
  AND2_X1 U186 ( .A1(n251), .A2(n303), .ZN(n298) );
  AOI21_X1 U187 ( .B1(net487913), .B2(n622), .A(n616), .ZN(n144) );
  NAND2_X1 U188 ( .A1(n433), .A2(n434), .ZN(n395) );
  NAND2_X1 U189 ( .A1(n441), .A2(n442), .ZN(n439) );
  NAND2_X1 U190 ( .A1(n325), .A2(n326), .ZN(n324) );
  INV_X1 U191 ( .A(n25), .ZN(n609) );
  NAND2_X1 U192 ( .A1(n13), .A2(n64), .ZN(n152) );
  NAND2_X1 U193 ( .A1(n352), .A2(n353), .ZN(n373) );
  AND3_X1 U194 ( .A1(net487908), .A2(n580), .A3(net487910), .ZN(net487907) );
  NAND2_X1 U195 ( .A1(n680), .A2(n653), .ZN(n406) );
  NAND2_X1 U196 ( .A1(n624), .A2(n681), .ZN(n181) );
  NAND2_X1 U197 ( .A1(n256), .A2(n257), .ZN(n300) );
  NAND2_X1 U198 ( .A1(n55), .A2(n167), .ZN(n154) );
  NAND2_X1 U199 ( .A1(n198), .A2(n185), .ZN(n188) );
  INV_X1 U200 ( .A(net487938), .ZN(n622) );
  NAND2_X1 U201 ( .A1(n291), .A2(n254), .ZN(n313) );
  NAND2_X1 U202 ( .A1(n286), .A2(n287), .ZN(n279) );
  NOR2_X1 U203 ( .A1(n293), .A2(n638), .ZN(n288) );
  INV_X1 U204 ( .A(n421), .ZN(n654) );
  XNOR2_X1 U205 ( .A(n446), .B(n445), .ZN(SUM[27]) );
  NAND2_X1 U206 ( .A1(n447), .A2(n436), .ZN(n446) );
  INV_X1 U207 ( .A(n360), .ZN(n650) );
  NAND2_X1 U208 ( .A1(n209), .A2(n168), .ZN(n208) );
  NOR2_X1 U209 ( .A1(n615), .A2(n617), .ZN(net487908) );
  INV_X1 U210 ( .A(net487913), .ZN(n617) );
  NAND2_X1 U211 ( .A1(n265), .A2(n266), .ZN(n264) );
  AOI21_X1 U212 ( .B1(n165), .B2(n166), .A(n569), .ZN(n163) );
  NAND2_X1 U213 ( .A1(n444), .A2(n443), .ZN(n453) );
  INV_X1 U214 ( .A(n303), .ZN(n637) );
  NAND2_X1 U215 ( .A1(n65), .A2(n9), .ZN(n74) );
  NOR2_X1 U216 ( .A1(n598), .A2(net487933), .ZN(n10) );
  INV_X1 U217 ( .A(net487940), .ZN(n598) );
  INV_X1 U218 ( .A(net487964), .ZN(n623) );
  NAND2_X1 U219 ( .A1(n162), .A2(net487998), .ZN(n161) );
  AND2_X1 U220 ( .A1(n268), .A2(n267), .ZN(n330) );
  INV_X1 U221 ( .A(n359), .ZN(n629) );
  INV_X1 U222 ( .A(n127), .ZN(n618) );
  INV_X1 U223 ( .A(n209), .ZN(n606) );
  INV_X1 U224 ( .A(n245), .ZN(n645) );
  NAND2_X1 U225 ( .A1(n406), .A2(n417), .ZN(n419) );
  NAND2_X1 U226 ( .A1(n279), .A2(n245), .ZN(n278) );
  INV_X1 U227 ( .A(n168), .ZN(n627) );
  AND2_X1 U228 ( .A1(n265), .A2(n266), .ZN(n26) );
  OAI21_X1 U229 ( .B1(n393), .B2(n394), .A(n395), .ZN(n389) );
  NAND2_X1 U230 ( .A1(n680), .A2(n653), .ZN(n388) );
  AND3_X1 U231 ( .A1(n392), .A2(n412), .A3(n421), .ZN(n390) );
  INV_X1 U232 ( .A(n254), .ZN(n638) );
  NAND2_X1 U233 ( .A1(n52), .A2(n53), .ZN(n143) );
  NOR2_X1 U234 ( .A1(n597), .A2(n147), .ZN(n53) );
  AND2_X1 U235 ( .A1(net487913), .A2(net487964), .ZN(n52) );
  INV_X1 U236 ( .A(n146), .ZN(n597) );
  INV_X1 U237 ( .A(n130), .ZN(n621) );
  INV_X1 U238 ( .A(n326), .ZN(n649) );
  INV_X1 U239 ( .A(n325), .ZN(n632) );
  NOR2_X1 U240 ( .A1(n605), .A2(n373), .ZN(n350) );
  INV_X1 U241 ( .A(n238), .ZN(n605) );
  AND2_X1 U242 ( .A1(n198), .A2(n207), .ZN(n14) );
  INV_X1 U243 ( .A(n157), .ZN(n610) );
  XNOR2_X1 U244 ( .A(n529), .B(n530), .ZN(SUM[15]) );
  NAND2_X1 U245 ( .A1(n531), .A2(n514), .ZN(n530) );
  NAND2_X1 U246 ( .A1(n510), .A2(n516), .ZN(n529) );
  NAND2_X1 U247 ( .A1(n515), .A2(n532), .ZN(n531) );
  XNOR2_X1 U248 ( .A(n503), .B(n402), .ZN(SUM[16]) );
  NAND2_X1 U249 ( .A1(n490), .A2(n487), .ZN(n503) );
  XNOR2_X1 U250 ( .A(n494), .B(n495), .ZN(SUM[19]) );
  NAND2_X1 U251 ( .A1(n489), .A2(n496), .ZN(n495) );
  NAND2_X1 U252 ( .A1(n484), .A2(n482), .ZN(n494) );
  NAND2_X1 U253 ( .A1(n483), .A2(n497), .ZN(n496) );
  XNOR2_X1 U254 ( .A(n470), .B(n469), .ZN(SUM[22]) );
  NAND2_X1 U255 ( .A1(n462), .A2(n459), .ZN(n470) );
  XNOR2_X1 U256 ( .A(n498), .B(n497), .ZN(SUM[18]) );
  NAND2_X1 U257 ( .A1(n483), .A2(n489), .ZN(n498) );
  XNOR2_X1 U258 ( .A(n499), .B(n500), .ZN(SUM[17]) );
  NOR2_X1 U259 ( .A1(n667), .A2(n666), .ZN(n500) );
  INV_X1 U260 ( .A(n488), .ZN(n667) );
  XNOR2_X1 U261 ( .A(n466), .B(n467), .ZN(SUM[23]) );
  NAND2_X1 U262 ( .A1(n459), .A2(n468), .ZN(n467) );
  NAND2_X1 U263 ( .A1(n462), .A2(n469), .ZN(n468) );
  INV_X1 U264 ( .A(n491), .ZN(n666) );
  XNOR2_X1 U265 ( .A(n533), .B(n532), .ZN(SUM[14]) );
  NAND2_X1 U266 ( .A1(n515), .A2(n514), .ZN(n533) );
  XNOR2_X1 U267 ( .A(n536), .B(n535), .ZN(SUM[13]) );
  NAND2_X1 U268 ( .A1(n520), .A2(n513), .ZN(n536) );
  XNOR2_X1 U269 ( .A(n477), .B(n476), .ZN(SUM[20]) );
  NAND2_X1 U270 ( .A1(n465), .A2(n464), .ZN(n477) );
  XNOR2_X1 U271 ( .A(n92), .B(n93), .ZN(SUM[7]) );
  NAND2_X1 U272 ( .A1(n96), .A2(n97), .ZN(n92) );
  NAND2_X1 U273 ( .A1(n94), .A2(n95), .ZN(n93) );
  NAND2_X1 U274 ( .A1(n98), .A2(n99), .ZN(n97) );
  XNOR2_X1 U275 ( .A(n333), .B(n334), .ZN(SUM[3]) );
  NAND2_X1 U276 ( .A1(n337), .A2(n338), .ZN(n333) );
  NAND2_X1 U277 ( .A1(n335), .A2(n336), .ZN(n334) );
  NAND2_X1 U278 ( .A1(n339), .A2(n340), .ZN(n338) );
  XNOR2_X1 U279 ( .A(n548), .B(n549), .ZN(SUM[11]) );
  NAND2_X1 U280 ( .A1(n544), .A2(n550), .ZN(n549) );
  NAND2_X1 U281 ( .A1(n545), .A2(n541), .ZN(n548) );
  NAND2_X1 U282 ( .A1(n547), .A2(n551), .ZN(n550) );
  XNOR2_X1 U283 ( .A(n492), .B(n686), .ZN(SUM[1]) );
  NAND2_X1 U284 ( .A1(n426), .A2(n425), .ZN(n492) );
  XNOR2_X1 U285 ( .A(n539), .B(n538), .ZN(SUM[12]) );
  NAND2_X1 U286 ( .A1(n519), .A2(n512), .ZN(n539) );
  XNOR2_X1 U287 ( .A(n88), .B(n89), .ZN(SUM[8]) );
  NAND2_X1 U288 ( .A1(n90), .A2(n91), .ZN(n88) );
  XNOR2_X1 U289 ( .A(n84), .B(n85), .ZN(SUM[9]) );
  NAND2_X1 U290 ( .A1(n86), .A2(n87), .ZN(n84) );
  XNOR2_X1 U291 ( .A(n137), .B(n105), .ZN(SUM[5]) );
  NAND2_X1 U292 ( .A1(n104), .A2(n103), .ZN(n137) );
  XNOR2_X1 U293 ( .A(n100), .B(n98), .ZN(SUM[6]) );
  NAND2_X1 U294 ( .A1(n99), .A2(n96), .ZN(n100) );
  XNOR2_X1 U295 ( .A(n552), .B(n551), .ZN(SUM[10]) );
  NAND2_X1 U296 ( .A1(n547), .A2(n544), .ZN(n552) );
  XNOR2_X1 U297 ( .A(n423), .B(n339), .ZN(SUM[2]) );
  NAND2_X1 U298 ( .A1(n340), .A2(n337), .ZN(n423) );
  XNOR2_X1 U299 ( .A(n214), .B(n527), .ZN(SUM[4]) );
  NAND2_X1 U300 ( .A1(n140), .A2(n139), .ZN(n214) );
  OAI21_X1 U301 ( .B1(n504), .B2(n505), .A(n506), .ZN(n402) );
  NOR2_X1 U302 ( .A1(n521), .A2(n673), .ZN(n504) );
  NAND4_X1 U303 ( .A1(n519), .A2(n520), .A3(n515), .A4(n516), .ZN(n505) );
  AOI21_X1 U304 ( .B1(n507), .B2(n508), .A(n669), .ZN(n506) );
  OAI21_X1 U305 ( .B1(n562), .B2(n563), .A(n336), .ZN(n527) );
  NAND2_X1 U306 ( .A1(n340), .A2(n335), .ZN(n563) );
  NOR2_X1 U307 ( .A1(n564), .A2(n565), .ZN(n562) );
  NAND2_X1 U308 ( .A1(n337), .A2(n425), .ZN(n565) );
  OAI21_X1 U309 ( .B1(n675), .B2(n674), .A(n87), .ZN(n551) );
  INV_X1 U310 ( .A(n85), .ZN(n675) );
  INV_X1 U311 ( .A(n86), .ZN(n674) );
  OAI21_X1 U312 ( .B1(n671), .B2(n670), .A(n513), .ZN(n532) );
  INV_X1 U313 ( .A(n535), .ZN(n671) );
  OAI21_X1 U314 ( .B1(n660), .B2(n659), .A(n463), .ZN(n469) );
  INV_X1 U315 ( .A(n460), .ZN(n659) );
  INV_X1 U316 ( .A(n473), .ZN(n660) );
  OAI21_X1 U317 ( .B1(n499), .B2(n666), .A(n488), .ZN(n497) );
  OAI21_X1 U318 ( .B1(n661), .B2(n662), .A(n464), .ZN(n473) );
  INV_X1 U319 ( .A(n465), .ZN(n661) );
  OAI21_X1 U320 ( .B1(n679), .B2(n684), .A(n139), .ZN(n105) );
  INV_X1 U321 ( .A(n140), .ZN(n679) );
  OAI21_X1 U322 ( .B1(n678), .B2(n677), .A(n103), .ZN(n98) );
  INV_X1 U323 ( .A(n105), .ZN(n678) );
  INV_X1 U324 ( .A(n104), .ZN(n677) );
  OAI21_X1 U325 ( .B1(n665), .B2(n481), .A(n482), .ZN(n397) );
  INV_X1 U326 ( .A(n485), .ZN(n665) );
  NAND2_X1 U327 ( .A1(n483), .A2(n484), .ZN(n481) );
  OAI211_X1 U328 ( .C1(n666), .C2(n487), .A(n488), .B(n489), .ZN(n485) );
  OAI21_X1 U329 ( .B1(n556), .B2(n557), .A(n94), .ZN(n525) );
  NAND2_X1 U330 ( .A1(n95), .A2(n96), .ZN(n557) );
  NOR2_X1 U331 ( .A1(n18), .A2(n558), .ZN(n556) );
  AND2_X1 U332 ( .A1(n103), .A2(n139), .ZN(n18) );
  NAND4_X1 U333 ( .A1(n140), .A2(n104), .A3(n99), .A4(n94), .ZN(n528) );
  NAND4_X1 U334 ( .A1(n490), .A2(n491), .A3(n483), .A4(n484), .ZN(n411) );
  NAND4_X1 U335 ( .A1(n465), .A2(n460), .A3(n462), .A4(n457), .ZN(n413) );
  NAND4_X1 U336 ( .A1(n392), .A2(n402), .A3(n403), .A4(n404), .ZN(n378) );
  NOR2_X1 U337 ( .A1(n407), .A2(n408), .ZN(n403) );
  NOR2_X1 U338 ( .A1(n652), .A2(n654), .ZN(n404) );
  NAND2_X1 U339 ( .A1(n664), .A2(n603), .ZN(n408) );
  NAND4_X1 U340 ( .A1(n86), .A2(n90), .A3(n547), .A4(n541), .ZN(n526) );
  AOI21_X1 U341 ( .B1(n109), .B2(n110), .A(n111), .ZN(n106) );
  NAND2_X1 U342 ( .A1(n112), .A2(n113), .ZN(n111) );
  OAI211_X1 U343 ( .C1(n670), .C2(n512), .A(n513), .B(n514), .ZN(n508) );
  NOR2_X1 U344 ( .A1(n685), .A2(n493), .ZN(n564) );
  INV_X1 U345 ( .A(n426), .ZN(n685) );
  NAND2_X1 U346 ( .A1(n555), .A2(n91), .ZN(n85) );
  NAND2_X1 U347 ( .A1(n89), .A2(n90), .ZN(n555) );
  NAND2_X1 U348 ( .A1(n537), .A2(n512), .ZN(n535) );
  NAND2_X1 U349 ( .A1(n538), .A2(n519), .ZN(n537) );
  NAND2_X1 U350 ( .A1(n424), .A2(n425), .ZN(n339) );
  NAND2_X1 U351 ( .A1(n426), .A2(n686), .ZN(n424) );
  NAND2_X1 U352 ( .A1(n541), .A2(n542), .ZN(n523) );
  NAND2_X1 U353 ( .A1(n87), .A2(n91), .ZN(n546) );
  INV_X1 U354 ( .A(n493), .ZN(n686) );
  AND2_X1 U355 ( .A1(n502), .A2(n487), .ZN(n499) );
  NAND2_X1 U356 ( .A1(n402), .A2(n490), .ZN(n502) );
  INV_X1 U357 ( .A(n520), .ZN(n670) );
  NAND2_X1 U358 ( .A1(n104), .A2(n99), .ZN(n558) );
  NAND2_X1 U359 ( .A1(n658), .A2(n412), .ZN(n407) );
  AND2_X1 U360 ( .A1(n516), .A2(n515), .ZN(n507) );
  INV_X1 U361 ( .A(n108), .ZN(n620) );
  INV_X1 U362 ( .A(n510), .ZN(n669) );
  INV_X1 U363 ( .A(n120), .ZN(n619) );
  OAI21_X1 U364 ( .B1(n82), .B2(n224), .A(n225), .ZN(n222) );
  AOI21_X1 U365 ( .B1(n287), .B2(n227), .A(n228), .ZN(n224) );
  NOR2_X1 U366 ( .A1(A[47]), .A2(B[47]), .ZN(n81) );
  NAND2_X1 U367 ( .A1(B[49]), .A2(A[49]), .ZN(n168) );
  NAND2_X1 U368 ( .A1(B[36]), .A2(A[36]), .ZN(n326) );
  NAND2_X1 U369 ( .A1(n356), .A2(n357), .ZN(n265) );
  AND2_X1 U371 ( .A1(n237), .A2(n361), .ZN(n356) );
  OAI211_X1 U372 ( .C1(n358), .C2(n359), .A(n360), .B(n368), .ZN(n357) );
  AOI21_X1 U373 ( .B1(n280), .B2(n281), .A(n83), .ZN(n277) );
  NAND2_X1 U374 ( .A1(B[24]), .A2(A[24]), .ZN(n442) );
  NAND2_X1 U375 ( .A1(A[47]), .A2(B[47]), .ZN(n223) );
  NAND2_X1 U376 ( .A1(n571), .A2(B[51]), .ZN(n180) );
  NAND2_X1 U377 ( .A1(A[50]), .A2(B[50]), .ZN(n205) );
  NAND2_X1 U378 ( .A1(B[48]), .A2(A[48]), .ZN(n209) );
  NAND2_X1 U380 ( .A1(B[40]), .A2(A[40]), .ZN(n257) );
  NAND2_X1 U381 ( .A1(A[34]), .A2(B[34]), .ZN(n368) );
  NAND4_X1 U382 ( .A1(n305), .A2(n291), .A3(n254), .A4(n262), .ZN(n233) );
  NAND2_X1 U383 ( .A1(B[32]), .A2(A[32]), .ZN(n359) );
  OR2_X1 U384 ( .A1(A[28]), .A2(B[28]), .ZN(n412) );
  NAND2_X1 U385 ( .A1(B[28]), .A2(A[28]), .ZN(n385) );
  OR2_X1 U386 ( .A1(B[21]), .A2(A[21]), .ZN(n460) );
  NAND2_X1 U387 ( .A1(B[25]), .A2(A[25]), .ZN(n441) );
  OR2_X1 U388 ( .A1(B[32]), .A2(A[32]), .ZN(n352) );
  NAND2_X1 U389 ( .A1(A[42]), .A2(B[42]), .ZN(n303) );
  NAND2_X1 U391 ( .A1(A[43]), .A2(B[43]), .ZN(n251) );
  NAND2_X1 U392 ( .A1(A[26]), .A2(B[26]), .ZN(n436) );
  OR2_X1 U393 ( .A1(A[47]), .A2(B[47]), .ZN(n16) );
  NAND2_X1 U394 ( .A1(B[52]), .A2(A[52]), .ZN(net487986) );
  NAND2_X1 U395 ( .A1(A[37]), .A2(B[37]), .ZN(n325) );
  NAND2_X1 U396 ( .A1(B[62]), .A2(A[62]), .ZN(n113) );
  NAND2_X1 U397 ( .A1(B[31]), .A2(A[31]), .ZN(n381) );
  NAND2_X1 U398 ( .A1(B[29]), .A2(A[29]), .ZN(n386) );
  OR2_X1 U399 ( .A1(A[31]), .A2(B[31]), .ZN(n392) );
  NAND2_X1 U400 ( .A1(A[38]), .A2(B[38]), .ZN(n328) );
  NAND2_X1 U401 ( .A1(B[22]), .A2(A[22]), .ZN(n459) );
  OR2_X1 U402 ( .A1(B[25]), .A2(A[25]), .ZN(n438) );
  OR2_X1 U403 ( .A1(A[23]), .A2(B[23]), .ZN(n457) );
  NAND2_X1 U404 ( .A1(B[55]), .A2(A[55]), .ZN(net487938) );
  OR2_X1 U405 ( .A1(B[49]), .A2(A[49]), .ZN(n185) );
  OR2_X1 U406 ( .A1(B[24]), .A2(A[24]), .ZN(n443) );
  OR2_X1 U407 ( .A1(B[29]), .A2(A[29]), .ZN(n421) );
  OR2_X1 U408 ( .A1(B[62]), .A2(A[62]), .ZN(n120) );
  OR2_X1 U409 ( .A1(B[50]), .A2(A[50]), .ZN(n169) );
  OR2_X1 U410 ( .A1(A[52]), .A2(B[52]), .ZN(n157) );
  OR2_X1 U411 ( .A1(B[35]), .A2(A[35]), .ZN(n238) );
  OR2_X1 U412 ( .A1(B[63]), .A2(A[63]), .ZN(n108) );
  NAND2_X1 U413 ( .A1(A[23]), .A2(B[23]), .ZN(n458) );
  OR2_X1 U414 ( .A1(A[27]), .A2(B[27]), .ZN(n433) );
  NAND2_X1 U415 ( .A1(B[39]), .A2(A[39]), .ZN(n327) );
  OR2_X1 U416 ( .A1(A[58]), .A2(B[58]), .ZN(n37) );
  OR2_X1 U417 ( .A1(B[60]), .A2(A[60]), .ZN(n130) );
  NAND2_X1 U418 ( .A1(n382), .A2(n383), .ZN(n380) );
  OAI211_X1 U419 ( .C1(n654), .C2(n385), .A(n386), .B(n387), .ZN(n383) );
  AND2_X1 U420 ( .A1(n392), .A2(n3), .ZN(n382) );
  INV_X1 U421 ( .A(n182), .ZN(n607) );
  NAND2_X1 U422 ( .A1(A[48]), .A2(B[48]), .ZN(n184) );
  INV_X1 U423 ( .A(n185), .ZN(n625) );
  OR2_X1 U424 ( .A1(A[43]), .A2(B[43]), .ZN(n72) );
  NOR2_X1 U425 ( .A1(A[46]), .A2(B[46]), .ZN(n596) );
  OR2_X1 U426 ( .A1(B[18]), .A2(A[18]), .ZN(n483) );
  OR2_X1 U427 ( .A1(B[14]), .A2(A[14]), .ZN(n515) );
  OR2_X1 U428 ( .A1(B[22]), .A2(A[22]), .ZN(n462) );
  OR2_X1 U429 ( .A1(B[19]), .A2(A[19]), .ZN(n484) );
  OR2_X1 U430 ( .A1(B[13]), .A2(A[13]), .ZN(n520) );
  OR2_X1 U431 ( .A1(B[16]), .A2(A[16]), .ZN(n490) );
  OR2_X1 U432 ( .A1(B[20]), .A2(A[20]), .ZN(n465) );
  OR2_X1 U433 ( .A1(B[15]), .A2(A[15]), .ZN(n516) );
  OR2_X1 U434 ( .A1(B[17]), .A2(A[17]), .ZN(n491) );
  OR2_X1 U435 ( .A1(B[6]), .A2(A[6]), .ZN(n99) );
  OR2_X1 U436 ( .A1(B[5]), .A2(A[5]), .ZN(n104) );
  OR2_X1 U437 ( .A1(B[10]), .A2(A[10]), .ZN(n547) );
  OR2_X1 U438 ( .A1(B[9]), .A2(A[9]), .ZN(n86) );
  OR2_X1 U439 ( .A1(B[11]), .A2(A[11]), .ZN(n541) );
  OR2_X1 U440 ( .A1(B[7]), .A2(A[7]), .ZN(n94) );
  OR2_X1 U441 ( .A1(B[8]), .A2(A[8]), .ZN(n90) );
  OR2_X1 U442 ( .A1(B[2]), .A2(A[2]), .ZN(n340) );
  OR2_X1 U443 ( .A1(B[12]), .A2(A[12]), .ZN(n519) );
  OR2_X1 U444 ( .A1(B[1]), .A2(A[1]), .ZN(n426) );
  OR2_X1 U445 ( .A1(B[4]), .A2(A[4]), .ZN(n140) );
  INV_X1 U446 ( .A(B[30]), .ZN(n680) );
  INV_X1 U447 ( .A(B[42]), .ZN(n683) );
  INV_X1 U448 ( .A(B[51]), .ZN(n681) );
  OR2_X1 U449 ( .A1(B[3]), .A2(A[3]), .ZN(n335) );
  INV_X1 U450 ( .A(B[46]), .ZN(n682) );
  OR2_X1 U451 ( .A1(B[0]), .A2(A[0]), .ZN(n560) );
  NAND2_X1 U452 ( .A1(B[1]), .A2(A[1]), .ZN(n425) );
  NAND2_X1 U453 ( .A1(B[8]), .A2(A[8]), .ZN(n91) );
  NAND2_X1 U454 ( .A1(B[12]), .A2(A[12]), .ZN(n512) );
  NAND2_X1 U455 ( .A1(B[14]), .A2(A[14]), .ZN(n514) );
  NAND2_X1 U456 ( .A1(B[20]), .A2(A[20]), .ZN(n464) );
  NAND2_X1 U457 ( .A1(B[13]), .A2(A[13]), .ZN(n513) );
  NAND2_X1 U458 ( .A1(B[6]), .A2(A[6]), .ZN(n96) );
  NAND2_X1 U459 ( .A1(B[17]), .A2(A[17]), .ZN(n488) );
  NAND2_X1 U460 ( .A1(B[18]), .A2(A[18]), .ZN(n489) );
  NAND2_X1 U461 ( .A1(B[21]), .A2(A[21]), .ZN(n463) );
  NAND2_X1 U462 ( .A1(B[9]), .A2(A[9]), .ZN(n87) );
  NAND2_X1 U463 ( .A1(B[2]), .A2(A[2]), .ZN(n337) );
  NAND2_X1 U464 ( .A1(B[0]), .A2(A[0]), .ZN(n493) );
  NAND2_X1 U465 ( .A1(B[16]), .A2(A[16]), .ZN(n487) );
  NAND2_X1 U466 ( .A1(B[4]), .A2(A[4]), .ZN(n139) );
  NAND2_X1 U467 ( .A1(B[5]), .A2(A[5]), .ZN(n103) );
  NAND2_X1 U468 ( .A1(B[10]), .A2(A[10]), .ZN(n544) );
  NAND2_X1 U469 ( .A1(B[3]), .A2(A[3]), .ZN(n336) );
  NAND2_X1 U470 ( .A1(B[19]), .A2(A[19]), .ZN(n482) );
  NAND2_X1 U471 ( .A1(B[7]), .A2(A[7]), .ZN(n95) );
  NAND2_X1 U472 ( .A1(B[15]), .A2(A[15]), .ZN(n510) );
  NAND2_X1 U473 ( .A1(B[11]), .A2(A[11]), .ZN(n545) );
  OAI21_X1 U474 ( .B1(n607), .B2(n179), .A(n180), .ZN(n177) );
  NAND2_X1 U475 ( .A1(B[54]), .A2(n568), .ZN(net487987) );
  OR2_X1 U476 ( .A1(B[33]), .A2(A[33]), .ZN(n353) );
  NOR2_X1 U477 ( .A1(A[33]), .A2(B[33]), .ZN(n358) );
  NAND2_X1 U478 ( .A1(B[33]), .A2(A[33]), .ZN(n360) );
  NAND2_X1 U479 ( .A1(B[30]), .A2(A[30]), .ZN(n417) );
  NAND2_X1 U480 ( .A1(B[30]), .A2(A[30]), .ZN(n387) );
  OR2_X1 U481 ( .A1(A[30]), .A2(B[30]), .ZN(n3) );
  INV_X1 U482 ( .A(A[30]), .ZN(n653) );
  OAI21_X1 U483 ( .B1(n601), .B2(n654), .A(n386), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n317), .A2(n270), .ZN(n258) );
  INV_X1 U485 ( .A(net487920), .ZN(n611) );
  XNOR2_X1 U486 ( .A(n211), .B(n210), .ZN(SUM[50]) );
  OAI21_X1 U487 ( .B1(n241), .B2(n242), .A(n243), .ZN(n220) );
  NAND2_X1 U488 ( .A1(n636), .A2(n683), .ZN(n262) );
  NAND2_X1 U489 ( .A1(n683), .A2(n636), .ZN(n252) );
  AOI21_X1 U490 ( .B1(n153), .B2(n154), .A(n569), .ZN(n151) );
  INV_X1 U491 ( .A(n169), .ZN(n628) );
  NAND2_X1 U492 ( .A1(n416), .A2(n417), .ZN(n415) );
  NAND2_X1 U493 ( .A1(B[63]), .A2(A[63]), .ZN(n112) );
  NOR2_X1 U494 ( .A1(B[53]), .A2(n570), .ZN(net487985) );
  NAND2_X1 U495 ( .A1(A[53]), .A2(B[53]), .ZN(net487988) );
  OR2_X1 U496 ( .A1(B[53]), .A2(A[53]), .ZN(n158) );
  OR2_X1 U497 ( .A1(A[53]), .A2(B[53]), .ZN(n174) );
  NOR2_X1 U498 ( .A1(n591), .A2(n611), .ZN(n141) );
  XNOR2_X1 U499 ( .A(n68), .B(n275), .ZN(SUM[46]) );
  INV_X1 U500 ( .A(A[42]), .ZN(n636) );
  XNOR2_X1 U501 ( .A(n295), .B(n60), .ZN(SUM[44]) );
  NAND2_X1 U502 ( .A1(n149), .A2(net487940), .ZN(n135) );
  XNOR2_X1 U503 ( .A(n135), .B(n148), .ZN(SUM[56]) );
  NAND2_X1 U504 ( .A1(n135), .A2(net487907), .ZN(n134) );
  XNOR2_X1 U505 ( .A(n575), .B(n349), .ZN(SUM[36]) );
  AND2_X1 U506 ( .A1(n270), .A2(n329), .ZN(n9) );
  NAND2_X1 U507 ( .A1(n329), .A2(n267), .ZN(n348) );
  XNOR2_X1 U508 ( .A(n203), .B(n202), .ZN(SUM[51]) );
  NAND4_X1 U509 ( .A1(n231), .A2(n229), .A3(n232), .A4(n46), .ZN(n221) );
  XNOR2_X1 U510 ( .A(n271), .B(n272), .ZN(SUM[47]) );
  INV_X1 U511 ( .A(n244), .ZN(n642) );
  NAND2_X1 U512 ( .A1(n253), .A2(n244), .ZN(n282) );
  NAND2_X1 U513 ( .A1(A[44]), .A2(B[44]), .ZN(n287) );
  AND3_X1 U514 ( .A1(n244), .A2(n72), .A3(n291), .ZN(n290) );
  NAND2_X1 U515 ( .A1(A[56]), .A2(B[56]), .ZN(net487918) );
  INV_X1 U516 ( .A(net487910), .ZN(n613) );
  INV_X1 U517 ( .A(n131), .ZN(n600) );
  INV_X1 U518 ( .A(n39), .ZN(n612) );
  OAI211_X1 U519 ( .C1(net487913), .C2(n614), .A(n37), .B(n578), .ZN(n34) );
  INV_X1 U520 ( .A(n578), .ZN(n615) );
  NAND2_X1 U521 ( .A1(net487921), .A2(net487913), .ZN(net487950) );
  NAND2_X1 U522 ( .A1(n120), .A2(n113), .ZN(n125) );
  NAND4_X1 U523 ( .A1(n267), .A2(n268), .A3(n576), .A4(n270), .ZN(n235) );
  NAND2_X1 U524 ( .A1(n268), .A2(n325), .ZN(n346) );
  NAND2_X1 U525 ( .A1(n268), .A2(n267), .ZN(n342) );
  AOI21_X1 U526 ( .B1(n649), .B2(n268), .A(n632), .ZN(n343) );
  NAND2_X1 U527 ( .A1(n205), .A2(n54), .ZN(n210) );
  OAI211_X1 U528 ( .C1(n625), .C2(n184), .A(n168), .B(n205), .ZN(n182) );
  AND2_X1 U529 ( .A1(n205), .A2(n168), .ZN(n55) );
  NAND2_X1 U530 ( .A1(net487983), .A2(net487984), .ZN(net487939) );
  XNOR2_X1 U531 ( .A(n125), .B(n124), .ZN(SUM[62]) );
  OAI211_X1 U532 ( .C1(n600), .C2(n621), .A(n116), .B(n117), .ZN(n110) );
  NAND2_X1 U533 ( .A1(n130), .A2(n117), .ZN(n132) );
  OAI21_X1 U534 ( .B1(n600), .B2(n621), .A(n117), .ZN(n128) );
  NAND2_X1 U535 ( .A1(B[60]), .A2(A[60]), .ZN(n117) );
  NOR2_X1 U536 ( .A1(n629), .A2(n230), .ZN(n372) );
  NAND4_X1 U537 ( .A1(n378), .A2(n379), .A3(n380), .A4(n381), .ZN(n230) );
  XNOR2_X1 U538 ( .A(n370), .B(n371), .ZN(SUM[34]) );
  OAI21_X1 U539 ( .B1(n372), .B2(n373), .A(n360), .ZN(n371) );
  AND2_X1 U540 ( .A1(A[46]), .A2(B[46]), .ZN(n82) );
  INV_X1 U541 ( .A(A[46]), .ZN(n648) );
  NAND2_X1 U542 ( .A1(net487981), .A2(net487987), .ZN(n170) );
  AND2_X1 U543 ( .A1(net487964), .A2(net487981), .ZN(net487983) );
  AND2_X1 U544 ( .A1(net487981), .A2(n174), .ZN(n162) );
  NOR2_X1 U545 ( .A1(n609), .A2(n152), .ZN(n190) );
  XNOR2_X1 U546 ( .A(n189), .B(n76), .ZN(SUM[53]) );
  XNOR2_X1 U547 ( .A(n318), .B(n321), .ZN(SUM[41]) );
  OAI21_X1 U548 ( .B1(n319), .B2(n320), .A(n257), .ZN(n318) );
  NAND2_X1 U549 ( .A1(n458), .A2(n457), .ZN(n466) );
  XNOR2_X1 U550 ( .A(n448), .B(n449), .ZN(SUM[26]) );
  NAND2_X1 U551 ( .A1(n581), .A2(n448), .ZN(n447) );
  NAND2_X1 U552 ( .A1(n458), .A2(n459), .ZN(n456) );
  AND2_X1 U553 ( .A1(A[45]), .A2(B[45]), .ZN(n83) );
  INV_X1 U554 ( .A(A[45]), .ZN(n644) );
  INV_X1 U555 ( .A(net487919), .ZN(n614) );
  NOR3_X1 U556 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n232) );
  INV_X1 U557 ( .A(n233), .ZN(n635) );
  NOR2_X1 U558 ( .A1(n81), .A2(n646), .ZN(n272) );
  NOR2_X1 U559 ( .A1(n596), .A2(n81), .ZN(n225) );
  NOR3_X1 U560 ( .A1(n81), .A2(n645), .A3(n642), .ZN(n231) );
  NAND2_X1 U561 ( .A1(A[57]), .A2(B[57]), .ZN(net487919) );
  AND2_X1 U562 ( .A1(net487988), .A2(n158), .ZN(n76) );
  OAI211_X1 U564 ( .C1(net487985), .C2(net487986), .A(net487988), .B(net487987), .ZN(net487984) );
  NAND2_X1 U565 ( .A1(net487988), .A2(net487986), .ZN(net487998) );
  NAND2_X1 U567 ( .A1(n437), .A2(n433), .ZN(n445) );
  XNOR2_X1 U568 ( .A(net487943), .B(n141), .ZN(SUM[58]) );
  XNOR2_X1 U569 ( .A(n283), .B(n284), .ZN(SUM[45]) );
  NOR2_X1 U570 ( .A1(n279), .A2(n285), .ZN(n283) );
  NAND2_X1 U571 ( .A1(n127), .A2(n116), .ZN(n129) );
  OR2_X1 U572 ( .A1(B[61]), .A2(A[61]), .ZN(n127) );
  AOI21_X1 U574 ( .B1(n62), .B2(n176), .A(n177), .ZN(n172) );
  AOI21_X1 U575 ( .B1(n274), .B2(n229), .A(n82), .ZN(n271) );
  OAI211_X1 U576 ( .C1(n615), .C2(net487918), .A(net487919), .B(net487920), 
        .ZN(net487915) );
  NAND2_X1 U583 ( .A1(net487913), .A2(net487918), .ZN(n148) );
  NAND2_X1 U584 ( .A1(net487918), .A2(net487938), .ZN(net487952) );
  INV_X1 U585 ( .A(net487918), .ZN(n616) );
  NOR2_X1 U586 ( .A1(n619), .A2(n618), .ZN(n109) );
  NAND2_X1 U588 ( .A1(n7), .A2(n120), .ZN(n123) );
  OAI21_X1 U590 ( .B1(n599), .B2(n618), .A(n116), .ZN(n7) );
  OAI21_X1 U591 ( .B1(n599), .B2(n618), .A(n116), .ZN(n124) );
  NAND2_X1 U592 ( .A1(A[58]), .A2(B[58]), .ZN(net487920) );
  AOI21_X1 U593 ( .B1(n198), .B2(n62), .A(n606), .ZN(n215) );
  OAI21_X1 U595 ( .B1(n172), .B2(n590), .A(n173), .ZN(n171) );
  NAND2_X1 U596 ( .A1(net487998), .A2(n158), .ZN(n173) );
  XNOR2_X1 U597 ( .A(n171), .B(n170), .ZN(SUM[54]) );
  AND2_X1 U598 ( .A1(n54), .A2(n175), .ZN(n64) );
  XNOR2_X1 U599 ( .A(n175), .B(n219), .ZN(SUM[48]) );
  NOR2_X1 U600 ( .A1(n191), .A2(n190), .ZN(n189) );
  OAI221_X1 U602 ( .B1(n610), .B2(n180), .C1(n193), .C2(n586), .A(net487986), 
        .ZN(n191) );
  AND2_X1 U603 ( .A1(n278), .A2(n277), .ZN(n68) );
  NAND2_X1 U604 ( .A1(n278), .A2(n277), .ZN(n274) );
  XNOR2_X1 U605 ( .A(net487930), .B(net487929), .ZN(SUM[59]) );
  NAND2_X1 U606 ( .A1(net487931), .A2(net487920), .ZN(net487930) );
  NAND2_X1 U608 ( .A1(A[27]), .A2(B[27]), .ZN(n437) );
  NOR2_X1 U610 ( .A1(n628), .A2(n71), .ZN(n165) );
  NOR2_X1 U611 ( .A1(n186), .A2(n71), .ZN(n176) );
  NOR2_X1 U612 ( .A1(n71), .A2(n628), .ZN(n153) );
  NOR2_X1 U613 ( .A1(n71), .A2(n188), .ZN(n13) );
  NOR2_X1 U614 ( .A1(n71), .A2(n188), .ZN(n70) );
  AND2_X1 U615 ( .A1(n26), .A2(n27), .ZN(n5) );
  NAND2_X1 U616 ( .A1(n26), .A2(n27), .ZN(n329) );
  NAND2_X1 U617 ( .A1(A[35]), .A2(B[35]), .ZN(n266) );
  OR2_X1 U619 ( .A1(A[35]), .A2(B[35]), .ZN(n361) );
  NAND4_X1 U620 ( .A1(n221), .A2(n220), .A3(n222), .A4(n223), .ZN(n61) );
  NAND4_X1 U621 ( .A1(n221), .A2(n220), .A3(n222), .A4(n223), .ZN(n62) );
  NAND4_X1 U622 ( .A1(n221), .A2(n222), .A3(n220), .A4(n223), .ZN(n175) );
  NOR2_X1 U624 ( .A1(net538236), .A2(net487952), .ZN(n142) );
  NAND2_X1 U625 ( .A1(net538236), .A2(net487913), .ZN(n145) );
  NOR2_X1 U626 ( .A1(n622), .A2(net538236), .ZN(n149) );
  XNOR2_X1 U627 ( .A(n308), .B(n309), .ZN(SUM[43]) );
  NAND2_X1 U628 ( .A1(n180), .A2(n181), .ZN(n202) );
  NAND2_X1 U629 ( .A1(n54), .A2(n181), .ZN(n179) );
  INV_X1 U630 ( .A(A[51]), .ZN(n624) );
  NAND2_X1 U631 ( .A1(B[41]), .A2(A[41]), .ZN(n256) );
  XNOR2_X1 U632 ( .A(n128), .B(n129), .ZN(SUM[61]) );
  INV_X1 U633 ( .A(n128), .ZN(n599) );
  NAND2_X1 U634 ( .A1(n133), .A2(n134), .ZN(n131) );
  NAND2_X1 U635 ( .A1(B[59]), .A2(A[59]), .ZN(n39) );
  NAND2_X1 U636 ( .A1(B[61]), .A2(A[61]), .ZN(n116) );
  NAND2_X1 U637 ( .A1(n648), .A2(n682), .ZN(n229) );
  NAND2_X1 U638 ( .A1(n682), .A2(n648), .ZN(n246) );
  XNOR2_X1 U639 ( .A(n215), .B(n216), .ZN(SUM[49]) );
  XNOR2_X1 U642 ( .A(n582), .B(n419), .ZN(SUM[30]) );
  XNOR2_X1 U643 ( .A(n422), .B(n428), .ZN(SUM[29]) );
  NAND2_X1 U644 ( .A1(n418), .A2(n406), .ZN(n416) );
  INV_X1 U645 ( .A(n422), .ZN(n601) );
  OR2_X1 U646 ( .A1(n10), .A2(n34), .ZN(net487931) );
  NAND2_X1 U647 ( .A1(n59), .A2(n151), .ZN(n146) );
  NOR2_X1 U648 ( .A1(n160), .A2(n159), .ZN(n78) );
  NAND2_X1 U649 ( .A1(n161), .A2(net487987), .ZN(n160) );
  XNOR2_X1 U650 ( .A(n78), .B(n79), .ZN(SUM[55]) );
  NOR2_X1 U651 ( .A1(net487948), .A2(n614), .ZN(net487943) );
  XNOR2_X1 U652 ( .A(n131), .B(n132), .ZN(SUM[60]) );
  AOI21_X1 U653 ( .B1(n136), .B2(net487915), .A(n612), .ZN(n133) );
  NOR2_X1 U654 ( .A1(n613), .A2(n591), .ZN(n136) );
endmodule


module RCA_NBIT64_5 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_5_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_4_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net447705, net447701, net447700, net447695, net447694, net447693,
         net447692, net447691, net447689, net447685, net447684, net447675,
         net447673, net447672, net447653, net447636, net447630, net537195,
         net537785, net447702, net447690, net447659, net447656, net535350,
         net447674, net447669, net447668, net447667, net447666, net447664,
         net447662, net447660, net447676, n1, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n17, n18, n19, n21, n23, n24, n28, n29, n30, n31, n32,
         n33, n40, n41, n42, n44, n45, n46, n47, n49, n51, n52, n54, n56, n57,
         n58, n60, n61, n62, n63, n64, n65, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n94, n95, n96, n97, n99, n100, n101, n102, n103, n106,
         n107, n108, n109, n111, n112, n113, n114, n116, n117, n118, n119,
         n120, n121, n122, n123, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n141, n142, n143, n144, n145,
         n146, n148, n149, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n163, n164, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n177, n178, n179, n182, n184, n186, n187, n188, n189,
         n190, n192, n193, n194, n195, n196, n199, n200, n201, n202, n203,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n223, n224, n225, n227, n228, n229, n230, n232,
         n233, n234, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n253, n254, n256, n258, n260,
         n263, n264, n265, n266, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n288, n289, n292, n297, n298, n300, n301, n302, n303, n304, n305,
         n306, n307, n310, n311, n312, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n335, n337, n338, n339, n342, n343, n344, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n358, n359, n360,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n378, n379, n381, n382, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n403, n405, n406, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n430, n431, n432, n433, n434, n435,
         n436, n437, n439, n441, n442, n443, n444, n445, n448, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n484, n485, n486, n487,
         n490, n491, n492, n493, n494, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  NAND3_X1 U11 ( .A1(n175), .A2(n174), .A3(n5), .ZN(n58) );
  NAND3_X1 U57 ( .A1(n241), .A2(n209), .A3(n210), .ZN(n234) );
  NAND3_X1 U87 ( .A1(n8), .A2(net537195), .A3(n9), .ZN(n30) );
  OR2_X2 U99 ( .A1(A[46]), .A2(B[46]), .ZN(n208) );
  OR2_X2 U101 ( .A1(A[53]), .A2(B[53]), .ZN(n123) );
  NAND3_X1 U130 ( .A1(n9), .A2(n8), .A3(net537195), .ZN(n118) );
  XOR2_X1 U246 ( .A(n107), .B(n108), .Z(SUM[63]) );
  XOR2_X1 U351 ( .A(n228), .B(n229), .Z(SUM[47]) );
  OR2_X2 U375 ( .A1(A[48]), .A2(B[48]), .ZN(n159) );
  OR2_X2 U382 ( .A1(A[49]), .A2(B[49]), .ZN(n160) );
  NAND3_X1 U520 ( .A1(n175), .A2(n171), .A3(n49), .ZN(n173) );
  NAND3_X1 U525 ( .A1(n184), .A2(n174), .A3(n175), .ZN(n182) );
  NAND3_X1 U527 ( .A1(n190), .A2(n189), .A3(n227), .ZN(n188) );
  NAND3_X1 U533 ( .A1(n224), .A2(n71), .A3(n52), .ZN(n216) );
  NAND3_X1 U537 ( .A1(n234), .A2(n207), .A3(n220), .ZN(n233) );
  NAND3_X1 U549 ( .A1(n270), .A2(n271), .A3(n224), .ZN(n269) );
  NAND3_X1 U591 ( .A1(n472), .A2(n473), .A3(n474), .ZN(n471) );
  NAND3_X1 U592 ( .A1(n475), .A2(n77), .A3(n476), .ZN(n472) );
  NAND3_X1 U597 ( .A1(n486), .A2(n87), .A3(n86), .ZN(n485) );
  NAND3_X1 U598 ( .A1(n95), .A2(n487), .A3(n90), .ZN(n486) );
  OR2_X2 U2 ( .A1(B[56]), .A2(A[56]), .ZN(net447673) );
  OR2_X2 U138 ( .A1(A[45]), .A2(B[45]), .ZN(n220) );
  CLKBUF_X1 U3 ( .A(A[31]), .Z(n497) );
  CLKBUF_X1 U4 ( .A(n62), .Z(n498) );
  INV_X1 U5 ( .A(n511), .ZN(n207) );
  NAND3_X1 U6 ( .A1(n219), .A2(n218), .A3(n500), .ZN(n175) );
  INV_X1 U7 ( .A(n276), .ZN(n556) );
  AND2_X1 U8 ( .A1(n490), .A2(n423), .ZN(SUM[0]) );
  BUF_X1 U9 ( .A(A[46]), .Z(n499) );
  AND2_X1 U10 ( .A1(n505), .A2(n217), .ZN(n500) );
  BUF_X1 U12 ( .A(A[47]), .Z(n506) );
  AND2_X1 U13 ( .A1(net447674), .A2(net447673), .ZN(n501) );
  OAI211_X1 U14 ( .C1(n529), .C2(n163), .A(n171), .B(n164), .ZN(n502) );
  AND2_X1 U15 ( .A1(A[54]), .A2(B[54]), .ZN(n503) );
  NOR2_X2 U16 ( .A1(B[41]), .A2(A[41]), .ZN(n61) );
  CLKBUF_X1 U17 ( .A(n552), .Z(n504) );
  AND4_X1 U18 ( .A1(n246), .A2(n245), .A3(n243), .A4(n244), .ZN(n505) );
  AND4_X1 U19 ( .A1(n246), .A2(n245), .A3(n243), .A4(n244), .ZN(n46) );
  NOR2_X1 U20 ( .A1(A[44]), .A2(B[44]), .ZN(n511) );
  OR2_X2 U21 ( .A1(B[37]), .A2(A[37]), .ZN(n270) );
  NAND3_X1 U22 ( .A1(n241), .A2(n209), .A3(n210), .ZN(n507) );
  OR2_X1 U23 ( .A1(A[57]), .A2(B[57]), .ZN(net447674) );
  OR2_X1 U24 ( .A1(A[52]), .A2(B[52]), .ZN(n120) );
  AND2_X1 U25 ( .A1(n187), .A2(n188), .ZN(n508) );
  OR2_X2 U26 ( .A1(A[40]), .A2(B[40]), .ZN(n243) );
  OR2_X1 U27 ( .A1(A[43]), .A2(B[43]), .ZN(n509) );
  OR2_X1 U28 ( .A1(A[43]), .A2(B[43]), .ZN(n246) );
  CLKBUF_X1 U29 ( .A(n21), .Z(n510) );
  OR2_X1 U30 ( .A1(B[54]), .A2(A[54]), .ZN(n119) );
  NOR2_X1 U31 ( .A1(B[54]), .A2(A[54]), .ZN(n47) );
  XNOR2_X1 U32 ( .A(n512), .B(net537195), .ZN(SUM[52]) );
  NAND2_X1 U33 ( .A1(n129), .A2(n120), .ZN(n512) );
  XNOR2_X1 U34 ( .A(n166), .B(n513), .ZN(SUM[51]) );
  NAND2_X1 U35 ( .A1(n157), .A2(n146), .ZN(n513) );
  OR2_X2 U36 ( .A1(A[50]), .A2(B[50]), .ZN(n158) );
  NAND3_X1 U37 ( .A1(net447676), .A2(n6), .A3(n501), .ZN(net447660) );
  INV_X1 U38 ( .A(n208), .ZN(n553) );
  AND2_X1 U39 ( .A1(net447673), .A2(net447674), .ZN(n514) );
  XNOR2_X1 U40 ( .A(n45), .B(n196), .ZN(SUM[48]) );
  XOR2_X1 U41 ( .A(n4), .B(n515), .Z(SUM[36]) );
  NOR2_X1 U42 ( .A1(n555), .A2(n556), .ZN(n515) );
  XOR2_X1 U43 ( .A(n230), .B(n516), .Z(SUM[46]) );
  NOR2_X1 U44 ( .A1(n73), .A2(n553), .ZN(n516) );
  INV_X1 U45 ( .A(n381), .ZN(n569) );
  INV_X1 U46 ( .A(n421), .ZN(n578) );
  OAI211_X1 U47 ( .C1(n200), .C2(n201), .A(n202), .B(n203), .ZN(n174) );
  OAI21_X1 U48 ( .B1(n569), .B2(n332), .A(n333), .ZN(n359) );
  NAND2_X1 U49 ( .A1(n44), .A2(n42), .ZN(net537195) );
  AOI21_X1 U50 ( .B1(n502), .B2(n143), .A(n525), .ZN(n44) );
  NAND2_X1 U51 ( .A1(n211), .A2(n263), .ZN(n242) );
  NOR2_X1 U52 ( .A1(n508), .A2(n178), .ZN(n184) );
  NAND2_X1 U53 ( .A1(n58), .A2(n31), .ZN(n42) );
  NOR2_X1 U54 ( .A1(n156), .A2(n155), .ZN(n31) );
  INV_X1 U55 ( .A(n378), .ZN(n566) );
  INV_X1 U56 ( .A(A[35]), .ZN(n565) );
  NAND2_X1 U58 ( .A1(n142), .A2(n152), .ZN(n121) );
  AOI21_X1 U59 ( .B1(n143), .B2(n144), .A(n525), .ZN(n152) );
  NAND2_X1 U60 ( .A1(n154), .A2(n58), .ZN(n142) );
  NOR2_X1 U61 ( .A1(n156), .A2(n155), .ZN(n154) );
  INV_X1 U62 ( .A(n170), .ZN(n530) );
  OAI21_X1 U63 ( .B1(n592), .B2(n457), .A(n454), .ZN(n80) );
  OAI21_X1 U64 ( .B1(n578), .B2(n344), .A(n574), .ZN(n395) );
  INV_X1 U65 ( .A(n335), .ZN(n574) );
  OAI21_X1 U66 ( .B1(n573), .B2(n338), .A(n337), .ZN(n381) );
  INV_X1 U67 ( .A(n395), .ZN(n573) );
  AOI21_X1 U68 ( .B1(n453), .B2(n454), .A(n455), .ZN(n448) );
  NAND2_X1 U69 ( .A1(n586), .A2(n456), .ZN(n453) );
  INV_X1 U70 ( .A(n457), .ZN(n586) );
  NAND2_X1 U71 ( .A1(n434), .A2(n435), .ZN(n421) );
  OAI21_X1 U72 ( .B1(n448), .B2(n583), .A(n10), .ZN(n434) );
  AOI21_X1 U73 ( .B1(n436), .B2(n437), .A(n579), .ZN(n435) );
  INV_X1 U74 ( .A(n452), .ZN(n583) );
  NAND2_X1 U75 ( .A1(n469), .A2(n452), .ZN(n467) );
  NAND2_X1 U76 ( .A1(n582), .A2(n80), .ZN(n469) );
  INV_X1 U77 ( .A(n455), .ZN(n582) );
  INV_X1 U78 ( .A(n456), .ZN(n592) );
  INV_X1 U79 ( .A(n338), .ZN(n568) );
  NOR2_X1 U80 ( .A1(n97), .A2(n540), .ZN(SUM[64]) );
  NOR2_X1 U81 ( .A1(n503), .A2(n47), .ZN(n138) );
  NOR2_X1 U82 ( .A1(n47), .A2(n136), .ZN(n133) );
  NOR2_X1 U83 ( .A1(n61), .A2(n549), .ZN(n260) );
  INV_X1 U84 ( .A(n250), .ZN(n549) );
  NAND2_X1 U85 ( .A1(n274), .A2(n224), .ZN(n65) );
  NAND2_X1 U86 ( .A1(n304), .A2(n301), .ZN(n314) );
  XOR2_X1 U88 ( .A(n33), .B(n292), .Z(SUM[37]) );
  NAND2_X1 U89 ( .A1(n328), .A2(n327), .ZN(n350) );
  NOR2_X1 U90 ( .A1(n526), .A2(n527), .ZN(n63) );
  INV_X1 U91 ( .A(n123), .ZN(n532) );
  NOR2_X1 U92 ( .A1(n537), .A2(net535350), .ZN(net447685) );
  NOR2_X1 U93 ( .A1(n533), .A2(n535), .ZN(n196) );
  XNOR2_X1 U94 ( .A(n237), .B(n238), .ZN(SUM[45]) );
  NOR2_X1 U95 ( .A1(n551), .A2(n504), .ZN(n238) );
  INV_X1 U96 ( .A(n220), .ZN(n551) );
  INV_X1 U97 ( .A(n103), .ZN(n539) );
  INV_X1 U98 ( .A(net537785), .ZN(n522) );
  INV_X1 U100 ( .A(n270), .ZN(n557) );
  OAI211_X1 U102 ( .C1(n70), .C2(n223), .A(n214), .B(n215), .ZN(n4) );
  NAND2_X1 U103 ( .A1(net447674), .A2(net447668), .ZN(net447700) );
  NOR2_X1 U104 ( .A1(n561), .A2(n560), .ZN(n254) );
  INV_X1 U105 ( .A(n509), .ZN(n560) );
  NAND4_X1 U106 ( .A1(n305), .A2(n304), .A3(n306), .A4(n307), .ZN(n223) );
  OAI21_X1 U107 ( .B1(n362), .B2(n12), .A(n363), .ZN(n333) );
  AND3_X1 U108 ( .A1(n366), .A2(n367), .A3(n368), .ZN(n12) );
  NAND2_X1 U109 ( .A1(n364), .A2(n365), .ZN(n362) );
  NAND2_X1 U110 ( .A1(n369), .A2(n370), .ZN(n367) );
  NOR2_X1 U111 ( .A1(n216), .A2(n223), .ZN(n217) );
  AND3_X1 U112 ( .A1(n208), .A2(n221), .A3(n220), .ZN(n219) );
  NAND2_X1 U113 ( .A1(n590), .A2(n554), .ZN(n218) );
  AOI21_X1 U114 ( .B1(n211), .B2(n212), .A(n548), .ZN(n200) );
  OR2_X1 U115 ( .A1(n216), .A2(n72), .ZN(n212) );
  INV_X1 U116 ( .A(n505), .ZN(n548) );
  AND2_X1 U117 ( .A1(n214), .A2(n215), .ZN(n72) );
  XNOR2_X1 U118 ( .A(n317), .B(n305), .ZN(SUM[32]) );
  NAND2_X1 U119 ( .A1(n306), .A2(n300), .ZN(n317) );
  XNOR2_X1 U120 ( .A(n310), .B(n311), .ZN(SUM[35]) );
  NAND2_X1 U121 ( .A1(n215), .A2(n303), .ZN(n311) );
  NAND2_X1 U122 ( .A1(n312), .A2(n301), .ZN(n310) );
  XOR2_X1 U123 ( .A(n517), .B(n351), .Z(SUM[29]) );
  NAND2_X1 U124 ( .A1(n326), .A2(n343), .ZN(n517) );
  XNOR2_X1 U125 ( .A(n347), .B(n346), .ZN(SUM[31]) );
  NAND2_X1 U126 ( .A1(n41), .A2(n321), .ZN(n346) );
  NAND2_X1 U127 ( .A1(n348), .A2(n327), .ZN(n347) );
  XNOR2_X1 U128 ( .A(n360), .B(n359), .ZN(SUM[28]) );
  NAND2_X1 U129 ( .A1(n342), .A2(n325), .ZN(n360) );
  XNOR2_X1 U131 ( .A(n379), .B(n378), .ZN(SUM[25]) );
  NAND2_X1 U132 ( .A1(n366), .A2(n369), .ZN(n379) );
  XNOR2_X1 U133 ( .A(n17), .B(n316), .ZN(SUM[33]) );
  NAND2_X1 U134 ( .A1(n307), .A2(n302), .ZN(n316) );
  OAI21_X1 U135 ( .B1(n544), .B2(n510), .A(n300), .ZN(n17) );
  XNOR2_X1 U136 ( .A(n285), .B(n286), .ZN(SUM[39]) );
  NOR2_X1 U137 ( .A1(n546), .A2(n545), .ZN(n286) );
  INV_X1 U139 ( .A(n288), .ZN(n546) );
  AND2_X1 U140 ( .A1(n199), .A2(n186), .ZN(n5) );
  XNOR2_X1 U141 ( .A(n40), .B(n258), .ZN(SUM[42]) );
  NAND2_X1 U142 ( .A1(n245), .A2(n251), .ZN(n258) );
  XNOR2_X1 U143 ( .A(n242), .B(n56), .ZN(SUM[40]) );
  NAND2_X1 U144 ( .A1(n243), .A2(n249), .ZN(n56) );
  XNOR2_X1 U145 ( .A(n372), .B(n373), .ZN(SUM[27]) );
  NAND2_X1 U146 ( .A1(n365), .A2(n374), .ZN(n372) );
  NAND2_X1 U147 ( .A1(n363), .A2(n364), .ZN(n373) );
  NAND2_X1 U148 ( .A1(n368), .A2(n375), .ZN(n374) );
  OAI211_X1 U149 ( .C1(n564), .C2(n300), .A(n301), .B(n302), .ZN(n298) );
  AND2_X1 U150 ( .A1(n303), .A2(n304), .ZN(n297) );
  INV_X1 U151 ( .A(n307), .ZN(n564) );
  NAND2_X1 U152 ( .A1(n46), .A2(n242), .ZN(n241) );
  AOI21_X1 U153 ( .B1(n275), .B2(n276), .A(n555), .ZN(n33) );
  OAI21_X1 U154 ( .B1(n521), .B2(n542), .A(n28), .ZN(net447653) );
  NAND4_X1 U155 ( .A1(n225), .A2(n224), .A3(n71), .A4(n4), .ZN(n263) );
  AND2_X1 U156 ( .A1(n288), .A2(n274), .ZN(n2) );
  OAI21_X1 U157 ( .B1(n351), .B2(n523), .A(n326), .ZN(n349) );
  OAI21_X1 U158 ( .B1(n167), .B2(n168), .A(n164), .ZN(n166) );
  OAI21_X1 U159 ( .B1(n566), .B2(n13), .A(n369), .ZN(n375) );
  OAI21_X1 U160 ( .B1(n567), .B2(n569), .A(n370), .ZN(n378) );
  INV_X1 U161 ( .A(n371), .ZN(n567) );
  INV_X1 U162 ( .A(n243), .ZN(n559) );
  AOI21_X1 U163 ( .B1(n266), .B2(n265), .A(n558), .ZN(n264) );
  AND4_X1 U164 ( .A1(n321), .A2(n319), .A3(n320), .A4(n318), .ZN(n21) );
  OAI21_X1 U165 ( .B1(n47), .B2(n131), .A(n130), .ZN(n135) );
  NOR2_X1 U166 ( .A1(n172), .A2(n173), .ZN(n167) );
  INV_X1 U167 ( .A(n178), .ZN(n534) );
  XNOR2_X1 U168 ( .A(n401), .B(n403), .ZN(SUM[21]) );
  NOR2_X1 U169 ( .A1(n572), .A2(n571), .ZN(n403) );
  INV_X1 U170 ( .A(n392), .ZN(n572) );
  AND2_X1 U171 ( .A1(n591), .A2(n565), .ZN(n70) );
  NAND2_X1 U172 ( .A1(n7), .A2(n30), .ZN(net537785) );
  NAND2_X1 U173 ( .A1(n187), .A2(n188), .ZN(n199) );
  AND2_X1 U174 ( .A1(n358), .A2(n325), .ZN(n351) );
  NAND2_X1 U175 ( .A1(n359), .A2(n342), .ZN(n358) );
  NAND2_X1 U176 ( .A1(n266), .A2(n52), .ZN(n211) );
  INV_X1 U177 ( .A(n302), .ZN(n563) );
  OAI21_X1 U178 ( .B1(n21), .B2(n544), .A(n300), .ZN(n315) );
  NAND2_X1 U179 ( .A1(n187), .A2(n188), .ZN(n177) );
  AND2_X1 U180 ( .A1(n208), .A2(n32), .ZN(n187) );
  NAND2_X1 U181 ( .A1(n554), .A2(n590), .ZN(n203) );
  NAND2_X1 U182 ( .A1(n209), .A2(n210), .ZN(n201) );
  NOR2_X1 U183 ( .A1(n511), .A2(n70), .ZN(n221) );
  NAND2_X1 U184 ( .A1(n591), .A2(n565), .ZN(n303) );
  NAND2_X1 U185 ( .A1(n247), .A2(n248), .ZN(n209) );
  AND2_X1 U186 ( .A1(n509), .A2(n57), .ZN(n247) );
  OAI211_X1 U187 ( .C1(n61), .C2(n249), .A(n250), .B(n251), .ZN(n248) );
  XNOR2_X1 U188 ( .A(n1), .B(n376), .ZN(SUM[26]) );
  OAI21_X1 U189 ( .B1(n566), .B2(n13), .A(n369), .ZN(n1) );
  NAND2_X1 U190 ( .A1(n368), .A2(n365), .ZN(n376) );
  INV_X1 U191 ( .A(n390), .ZN(n571) );
  INV_X1 U192 ( .A(n29), .ZN(n542) );
  INV_X1 U193 ( .A(n146), .ZN(n525) );
  INV_X1 U194 ( .A(n306), .ZN(n544) );
  INV_X1 U195 ( .A(n273), .ZN(n555) );
  INV_X1 U196 ( .A(n343), .ZN(n523) );
  AND2_X1 U197 ( .A1(n276), .A2(n270), .ZN(n71) );
  INV_X1 U198 ( .A(n131), .ZN(n531) );
  NAND2_X1 U199 ( .A1(n120), .A2(n123), .ZN(n136) );
  NAND2_X1 U200 ( .A1(n69), .A2(n330), .ZN(n319) );
  OAI21_X1 U201 ( .B1(n331), .B2(n332), .A(n333), .ZN(n330) );
  AOI21_X1 U202 ( .B1(n568), .B2(n335), .A(n570), .ZN(n331) );
  INV_X1 U203 ( .A(n337), .ZN(n570) );
  INV_X1 U204 ( .A(n112), .ZN(n541) );
  INV_X1 U205 ( .A(n164), .ZN(n526) );
  NAND2_X1 U206 ( .A1(n170), .A2(n171), .ZN(n169) );
  AND2_X1 U207 ( .A1(n119), .A2(n120), .ZN(n9) );
  INV_X1 U208 ( .A(n239), .ZN(n550) );
  INV_X1 U209 ( .A(n210), .ZN(n561) );
  AND2_X1 U210 ( .A1(n225), .A2(n243), .ZN(n265) );
  INV_X1 U211 ( .A(n249), .ZN(n558) );
  NAND2_X1 U212 ( .A1(n322), .A2(n323), .ZN(n320) );
  OAI211_X1 U213 ( .C1(n523), .C2(n325), .A(n326), .B(n327), .ZN(n323) );
  AND2_X1 U214 ( .A1(n41), .A2(n328), .ZN(n322) );
  INV_X1 U215 ( .A(n159), .ZN(n535) );
  INV_X1 U216 ( .A(n52), .ZN(n545) );
  INV_X1 U217 ( .A(n171), .ZN(n528) );
  AND2_X1 U218 ( .A1(n123), .A2(n120), .ZN(n60) );
  INV_X1 U219 ( .A(n251), .ZN(n562) );
  INV_X1 U220 ( .A(n274), .ZN(n547) );
  XNOR2_X1 U221 ( .A(n424), .B(n425), .ZN(SUM[19]) );
  NAND2_X1 U222 ( .A1(n415), .A2(n426), .ZN(n424) );
  NAND2_X1 U223 ( .A1(n410), .A2(n412), .ZN(n425) );
  NAND2_X1 U224 ( .A1(n427), .A2(n411), .ZN(n426) );
  XNOR2_X1 U225 ( .A(n458), .B(n459), .ZN(SUM[15]) );
  NAND2_X1 U226 ( .A1(n460), .A2(n443), .ZN(n459) );
  NAND2_X1 U227 ( .A1(n439), .A2(n445), .ZN(n458) );
  NAND2_X1 U228 ( .A1(n444), .A2(n461), .ZN(n460) );
  XNOR2_X1 U229 ( .A(n396), .B(n397), .ZN(SUM[23]) );
  NAND2_X1 U230 ( .A1(n388), .A2(n398), .ZN(n397) );
  NAND2_X1 U231 ( .A1(n387), .A2(n386), .ZN(n396) );
  NAND2_X1 U232 ( .A1(n391), .A2(n399), .ZN(n398) );
  XNOR2_X1 U233 ( .A(n431), .B(n430), .ZN(SUM[17]) );
  NAND2_X1 U234 ( .A1(n420), .A2(n416), .ZN(n431) );
  XNOR2_X1 U235 ( .A(n382), .B(n381), .ZN(SUM[24]) );
  NAND2_X1 U236 ( .A1(n371), .A2(n370), .ZN(n382) );
  XNOR2_X1 U237 ( .A(n462), .B(n461), .ZN(SUM[14]) );
  NAND2_X1 U238 ( .A1(n444), .A2(n443), .ZN(n462) );
  XNOR2_X1 U239 ( .A(n400), .B(n399), .ZN(SUM[22]) );
  NAND2_X1 U240 ( .A1(n391), .A2(n388), .ZN(n400) );
  XNOR2_X1 U241 ( .A(n433), .B(n421), .ZN(SUM[16]) );
  NAND2_X1 U242 ( .A1(n418), .A2(n419), .ZN(n433) );
  XNOR2_X1 U243 ( .A(n428), .B(n427), .ZN(SUM[18]) );
  NAND2_X1 U244 ( .A1(n411), .A2(n415), .ZN(n428) );
  XNOR2_X1 U245 ( .A(n465), .B(n464), .ZN(SUM[13]) );
  NAND2_X1 U247 ( .A1(n451), .A2(n442), .ZN(n465) );
  XNOR2_X1 U248 ( .A(n406), .B(n395), .ZN(SUM[20]) );
  NAND2_X1 U249 ( .A1(n394), .A2(n393), .ZN(n406) );
  XNOR2_X1 U250 ( .A(n83), .B(n84), .ZN(SUM[7]) );
  NAND2_X1 U251 ( .A1(n87), .A2(n88), .ZN(n83) );
  NAND2_X1 U252 ( .A1(n85), .A2(n86), .ZN(n84) );
  NAND2_X1 U253 ( .A1(n89), .A2(n90), .ZN(n88) );
  XNOR2_X1 U254 ( .A(n277), .B(n278), .ZN(SUM[3]) );
  NAND2_X1 U255 ( .A1(n281), .A2(n282), .ZN(n277) );
  NAND2_X1 U256 ( .A1(n279), .A2(n280), .ZN(n278) );
  NAND2_X1 U257 ( .A1(n283), .A2(n284), .ZN(n282) );
  XNOR2_X1 U258 ( .A(n477), .B(n478), .ZN(SUM[11]) );
  NAND2_X1 U259 ( .A1(n473), .A2(n479), .ZN(n478) );
  NAND2_X1 U260 ( .A1(n474), .A2(n470), .ZN(n477) );
  NAND2_X1 U261 ( .A1(n476), .A2(n480), .ZN(n479) );
  XNOR2_X1 U262 ( .A(n422), .B(n594), .ZN(SUM[1]) );
  NAND2_X1 U263 ( .A1(n355), .A2(n354), .ZN(n422) );
  XNOR2_X1 U264 ( .A(n468), .B(n467), .ZN(SUM[12]) );
  NAND2_X1 U265 ( .A1(n450), .A2(n441), .ZN(n468) );
  XNOR2_X1 U266 ( .A(n79), .B(n80), .ZN(SUM[8]) );
  NAND2_X1 U267 ( .A1(n81), .A2(n82), .ZN(n79) );
  XNOR2_X1 U268 ( .A(n114), .B(n96), .ZN(SUM[5]) );
  NAND2_X1 U269 ( .A1(n95), .A2(n94), .ZN(n114) );
  XNOR2_X1 U270 ( .A(n75), .B(n76), .ZN(SUM[9]) );
  NAND2_X1 U271 ( .A1(n77), .A2(n78), .ZN(n75) );
  XNOR2_X1 U272 ( .A(n91), .B(n89), .ZN(SUM[6]) );
  NAND2_X1 U273 ( .A1(n90), .A2(n87), .ZN(n91) );
  XNOR2_X1 U274 ( .A(n481), .B(n480), .ZN(SUM[10]) );
  NAND2_X1 U275 ( .A1(n476), .A2(n473), .ZN(n481) );
  XNOR2_X1 U276 ( .A(n352), .B(n283), .ZN(SUM[2]) );
  NAND2_X1 U277 ( .A1(n284), .A2(n281), .ZN(n352) );
  XNOR2_X1 U278 ( .A(n192), .B(n456), .ZN(SUM[4]) );
  NAND2_X1 U279 ( .A1(n117), .A2(n116), .ZN(n192) );
  OAI21_X1 U280 ( .B1(n491), .B2(n492), .A(n280), .ZN(n456) );
  NAND2_X1 U281 ( .A1(n284), .A2(n279), .ZN(n492) );
  NOR2_X1 U282 ( .A1(n493), .A2(n494), .ZN(n491) );
  NAND2_X1 U283 ( .A1(n281), .A2(n354), .ZN(n494) );
  OAI21_X1 U284 ( .B1(n585), .B2(n584), .A(n78), .ZN(n480) );
  INV_X1 U285 ( .A(n76), .ZN(n585) );
  INV_X1 U286 ( .A(n77), .ZN(n584) );
  OAI21_X1 U287 ( .B1(n581), .B2(n580), .A(n442), .ZN(n461) );
  INV_X1 U288 ( .A(n464), .ZN(n581) );
  OAI21_X1 U289 ( .B1(n401), .B2(n571), .A(n392), .ZN(n399) );
  OAI21_X1 U290 ( .B1(n589), .B2(n592), .A(n116), .ZN(n96) );
  INV_X1 U291 ( .A(n117), .ZN(n589) );
  OAI21_X1 U292 ( .B1(n588), .B2(n587), .A(n94), .ZN(n89) );
  INV_X1 U293 ( .A(n95), .ZN(n587) );
  INV_X1 U294 ( .A(n96), .ZN(n588) );
  OAI21_X1 U295 ( .B1(n577), .B2(n576), .A(n416), .ZN(n427) );
  INV_X1 U296 ( .A(n430), .ZN(n577) );
  NAND4_X1 U297 ( .A1(n394), .A2(n391), .A3(n390), .A4(n386), .ZN(n338) );
  NAND4_X1 U298 ( .A1(n371), .A2(n366), .A3(n368), .A4(n363), .ZN(n332) );
  OAI21_X1 U299 ( .B1(n408), .B2(n409), .A(n410), .ZN(n335) );
  NAND2_X1 U300 ( .A1(n411), .A2(n412), .ZN(n409) );
  NOR2_X1 U301 ( .A1(n413), .A2(n414), .ZN(n408) );
  NAND2_X1 U302 ( .A1(n415), .A2(n416), .ZN(n414) );
  OAI21_X1 U303 ( .B1(n384), .B2(n385), .A(n386), .ZN(n337) );
  NAND2_X1 U304 ( .A1(n387), .A2(n388), .ZN(n385) );
  NOR2_X1 U305 ( .A1(n11), .A2(n389), .ZN(n384) );
  AND2_X1 U306 ( .A1(n392), .A2(n393), .ZN(n11) );
  NAND4_X1 U307 ( .A1(n419), .A2(n420), .A3(n411), .A4(n412), .ZN(n344) );
  NAND4_X1 U308 ( .A1(n117), .A2(n95), .A3(n90), .A4(n85), .ZN(n457) );
  NAND4_X1 U309 ( .A1(n77), .A2(n81), .A3(n476), .A4(n470), .ZN(n455) );
  OAI211_X1 U310 ( .C1(n580), .C2(n441), .A(n442), .B(n443), .ZN(n437) );
  AOI21_X1 U311 ( .B1(n100), .B2(net447630), .A(n101), .ZN(n97) );
  NAND2_X1 U312 ( .A1(n102), .A2(n103), .ZN(n101) );
  NOR2_X1 U313 ( .A1(n538), .A2(n541), .ZN(n100) );
  OAI211_X1 U314 ( .C1(n521), .C2(n542), .A(net447636), .B(n28), .ZN(net447630) );
  NAND4_X1 U315 ( .A1(n339), .A2(n575), .A3(n524), .A4(n69), .ZN(n318) );
  INV_X1 U316 ( .A(n344), .ZN(n575) );
  INV_X1 U317 ( .A(n332), .ZN(n524) );
  NOR2_X1 U318 ( .A1(n578), .A2(n338), .ZN(n339) );
  NOR2_X1 U319 ( .A1(n576), .A2(n418), .ZN(n413) );
  NOR2_X1 U320 ( .A1(n593), .A2(n423), .ZN(n493) );
  INV_X1 U321 ( .A(n355), .ZN(n593) );
  NAND2_X1 U322 ( .A1(n484), .A2(n82), .ZN(n76) );
  NAND2_X1 U323 ( .A1(n80), .A2(n81), .ZN(n484) );
  NAND2_X1 U324 ( .A1(n466), .A2(n441), .ZN(n464) );
  NAND2_X1 U325 ( .A1(n467), .A2(n450), .ZN(n466) );
  NAND2_X1 U326 ( .A1(n432), .A2(n418), .ZN(n430) );
  NAND2_X1 U327 ( .A1(n421), .A2(n419), .ZN(n432) );
  NAND2_X1 U328 ( .A1(n353), .A2(n354), .ZN(n283) );
  NAND2_X1 U329 ( .A1(n355), .A2(n594), .ZN(n353) );
  NAND2_X1 U330 ( .A1(n470), .A2(n471), .ZN(n452) );
  NAND2_X1 U331 ( .A1(n78), .A2(n82), .ZN(n475) );
  NAND2_X1 U332 ( .A1(n85), .A2(n485), .ZN(n454) );
  NAND2_X1 U333 ( .A1(n94), .A2(n116), .ZN(n487) );
  INV_X1 U334 ( .A(n423), .ZN(n594) );
  AND2_X1 U335 ( .A1(n405), .A2(n393), .ZN(n401) );
  NAND2_X1 U336 ( .A1(n395), .A2(n394), .ZN(n405) );
  INV_X1 U337 ( .A(n420), .ZN(n576) );
  INV_X1 U338 ( .A(n451), .ZN(n580) );
  NAND2_X1 U339 ( .A1(n390), .A2(n391), .ZN(n389) );
  AND4_X1 U340 ( .A1(n450), .A2(n451), .A3(n444), .A4(n445), .ZN(n10) );
  AND2_X1 U341 ( .A1(n445), .A2(n444), .ZN(n436) );
  INV_X1 U342 ( .A(n99), .ZN(n540) );
  INV_X1 U343 ( .A(n439), .ZN(n579) );
  NAND2_X1 U344 ( .A1(n499), .A2(B[46]), .ZN(n227) );
  NOR2_X1 U345 ( .A1(A[25]), .A2(B[25]), .ZN(n13) );
  NAND2_X1 U346 ( .A1(B[25]), .A2(A[25]), .ZN(n369) );
  NAND2_X1 U347 ( .A1(B[32]), .A2(A[32]), .ZN(n300) );
  NAND2_X1 U348 ( .A1(A[49]), .A2(B[49]), .ZN(n171) );
  NAND2_X1 U349 ( .A1(B[41]), .A2(A[41]), .ZN(n250) );
  OR2_X1 U350 ( .A1(A[38]), .A2(B[38]), .ZN(n224) );
  NAND2_X1 U352 ( .A1(A[40]), .A2(B[40]), .ZN(n249) );
  NAND2_X1 U353 ( .A1(B[34]), .A2(A[34]), .ZN(n301) );
  OR2_X1 U354 ( .A1(B[33]), .A2(A[33]), .ZN(n307) );
  NAND2_X1 U355 ( .A1(B[35]), .A2(A[35]), .ZN(n215) );
  NAND2_X1 U356 ( .A1(B[30]), .A2(A[30]), .ZN(n327) );
  NAND2_X1 U357 ( .A1(B[42]), .A2(A[42]), .ZN(n251) );
  NAND2_X1 U358 ( .A1(B[24]), .A2(A[24]), .ZN(n370) );
  NAND2_X1 U359 ( .A1(B[26]), .A2(A[26]), .ZN(n365) );
  OR2_X1 U360 ( .A1(B[26]), .A2(A[26]), .ZN(n368) );
  NAND2_X1 U361 ( .A1(B[33]), .A2(A[33]), .ZN(n302) );
  NAND2_X1 U362 ( .A1(A[43]), .A2(B[43]), .ZN(n210) );
  NAND2_X1 U363 ( .A1(A[38]), .A2(B[38]), .ZN(n274) );
  NAND2_X1 U364 ( .A1(B[62]), .A2(A[62]), .ZN(n103) );
  OR2_X1 U365 ( .A1(A[34]), .A2(B[34]), .ZN(n304) );
  NAND2_X1 U366 ( .A1(B[51]), .A2(A[51]), .ZN(n146) );
  NAND2_X1 U367 ( .A1(B[28]), .A2(A[28]), .ZN(n325) );
  NAND2_X1 U368 ( .A1(B[29]), .A2(A[29]), .ZN(n326) );
  OR2_X1 U369 ( .A1(B[27]), .A2(A[27]), .ZN(n363) );
  OR2_X1 U370 ( .A1(B[32]), .A2(A[32]), .ZN(n306) );
  OR2_X1 U371 ( .A1(B[21]), .A2(A[21]), .ZN(n390) );
  NAND2_X1 U372 ( .A1(A[48]), .A2(B[48]), .ZN(n163) );
  NAND2_X1 U373 ( .A1(A[27]), .A2(B[27]), .ZN(n364) );
  OR2_X1 U374 ( .A1(B[30]), .A2(A[30]), .ZN(n328) );
  AND3_X1 U376 ( .A1(n329), .A2(n328), .A3(n51), .ZN(n69) );
  AND2_X1 U377 ( .A1(n343), .A2(n342), .ZN(n51) );
  OR2_X1 U378 ( .A1(B[36]), .A2(A[36]), .ZN(n276) );
  OR2_X1 U379 ( .A1(B[39]), .A2(A[39]), .ZN(n52) );
  NAND2_X1 U380 ( .A1(A[39]), .A2(B[39]), .ZN(n288) );
  OR2_X1 U381 ( .A1(B[41]), .A2(A[41]), .ZN(n244) );
  OR2_X1 U383 ( .A1(B[28]), .A2(A[28]), .ZN(n342) );
  OR2_X1 U384 ( .A1(A[25]), .A2(B[25]), .ZN(n366) );
  NOR2_X1 U385 ( .A1(A[57]), .A2(B[57]), .ZN(net447666) );
  NAND2_X1 U386 ( .A1(B[36]), .A2(A[36]), .ZN(n273) );
  OR2_X1 U387 ( .A1(A[29]), .A2(B[29]), .ZN(n343) );
  AND2_X1 U388 ( .A1(B[46]), .A2(n499), .ZN(n73) );
  OR2_X1 U389 ( .A1(A[51]), .A2(B[51]), .ZN(n157) );
  OR2_X1 U390 ( .A1(B[42]), .A2(A[42]), .ZN(n245) );
  OR2_X1 U391 ( .A1(B[62]), .A2(A[62]), .ZN(n106) );
  OR2_X1 U392 ( .A1(A[31]), .A2(B[31]), .ZN(n41) );
  OR2_X1 U393 ( .A1(B[63]), .A2(A[63]), .ZN(n99) );
  OR2_X1 U394 ( .A1(A[39]), .A2(B[39]), .ZN(n225) );
  OR2_X1 U395 ( .A1(B[42]), .A2(A[42]), .ZN(n57) );
  AND2_X1 U396 ( .A1(n122), .A2(n123), .ZN(n8) );
  OR2_X1 U397 ( .A1(B[18]), .A2(A[18]), .ZN(n411) );
  OR2_X1 U398 ( .A1(B[22]), .A2(A[22]), .ZN(n391) );
  OR2_X1 U399 ( .A1(B[14]), .A2(A[14]), .ZN(n444) );
  OR2_X1 U400 ( .A1(B[19]), .A2(A[19]), .ZN(n412) );
  OR2_X1 U401 ( .A1(B[23]), .A2(A[23]), .ZN(n386) );
  OR2_X1 U402 ( .A1(B[16]), .A2(A[16]), .ZN(n419) );
  OR2_X1 U403 ( .A1(B[13]), .A2(A[13]), .ZN(n451) );
  OR2_X1 U404 ( .A1(B[17]), .A2(A[17]), .ZN(n420) );
  OR2_X1 U405 ( .A1(B[20]), .A2(A[20]), .ZN(n394) );
  OR2_X1 U406 ( .A1(B[24]), .A2(A[24]), .ZN(n371) );
  OR2_X1 U407 ( .A1(B[15]), .A2(A[15]), .ZN(n445) );
  OR2_X1 U408 ( .A1(B[6]), .A2(A[6]), .ZN(n90) );
  OR2_X1 U409 ( .A1(B[10]), .A2(A[10]), .ZN(n476) );
  OR2_X1 U410 ( .A1(B[5]), .A2(A[5]), .ZN(n95) );
  OR2_X1 U411 ( .A1(B[9]), .A2(A[9]), .ZN(n77) );
  OR2_X1 U412 ( .A1(B[11]), .A2(A[11]), .ZN(n470) );
  OR2_X1 U413 ( .A1(B[7]), .A2(A[7]), .ZN(n85) );
  OR2_X1 U414 ( .A1(B[8]), .A2(A[8]), .ZN(n81) );
  OR2_X1 U415 ( .A1(B[2]), .A2(A[2]), .ZN(n284) );
  OR2_X1 U416 ( .A1(B[12]), .A2(A[12]), .ZN(n450) );
  OR2_X1 U417 ( .A1(B[1]), .A2(A[1]), .ZN(n355) );
  OR2_X1 U418 ( .A1(B[4]), .A2(A[4]), .ZN(n117) );
  INV_X1 U419 ( .A(B[47]), .ZN(n590) );
  INV_X1 U420 ( .A(B[35]), .ZN(n591) );
  OR2_X1 U421 ( .A1(B[3]), .A2(A[3]), .ZN(n279) );
  OR2_X1 U422 ( .A1(B[0]), .A2(A[0]), .ZN(n490) );
  NAND2_X1 U423 ( .A1(B[1]), .A2(A[1]), .ZN(n354) );
  NAND2_X1 U424 ( .A1(B[8]), .A2(A[8]), .ZN(n82) );
  NAND2_X1 U425 ( .A1(B[12]), .A2(A[12]), .ZN(n441) );
  NAND2_X1 U426 ( .A1(B[14]), .A2(A[14]), .ZN(n443) );
  NAND2_X1 U427 ( .A1(B[17]), .A2(A[17]), .ZN(n416) );
  NAND2_X1 U428 ( .A1(B[4]), .A2(A[4]), .ZN(n116) );
  NAND2_X1 U429 ( .A1(B[13]), .A2(A[13]), .ZN(n442) );
  NAND2_X1 U430 ( .A1(B[22]), .A2(A[22]), .ZN(n388) );
  NAND2_X1 U431 ( .A1(B[16]), .A2(A[16]), .ZN(n418) );
  NAND2_X1 U432 ( .A1(B[5]), .A2(A[5]), .ZN(n94) );
  NAND2_X1 U433 ( .A1(B[9]), .A2(A[9]), .ZN(n78) );
  NAND2_X1 U434 ( .A1(B[18]), .A2(A[18]), .ZN(n415) );
  NAND2_X1 U435 ( .A1(B[2]), .A2(A[2]), .ZN(n281) );
  NAND2_X1 U436 ( .A1(B[0]), .A2(A[0]), .ZN(n423) );
  NAND2_X1 U437 ( .A1(B[6]), .A2(A[6]), .ZN(n87) );
  NAND2_X1 U438 ( .A1(B[10]), .A2(A[10]), .ZN(n473) );
  NAND2_X1 U439 ( .A1(B[21]), .A2(A[21]), .ZN(n392) );
  NAND2_X1 U440 ( .A1(B[20]), .A2(A[20]), .ZN(n393) );
  NAND2_X1 U441 ( .A1(B[3]), .A2(A[3]), .ZN(n280) );
  NAND2_X1 U442 ( .A1(B[15]), .A2(A[15]), .ZN(n439) );
  NAND2_X1 U443 ( .A1(B[19]), .A2(A[19]), .ZN(n410) );
  NAND2_X1 U444 ( .A1(B[23]), .A2(A[23]), .ZN(n387) );
  NAND2_X1 U445 ( .A1(B[7]), .A2(A[7]), .ZN(n86) );
  NAND2_X1 U446 ( .A1(B[11]), .A2(A[11]), .ZN(n474) );
  NAND2_X1 U447 ( .A1(A[53]), .A2(B[53]), .ZN(n131) );
  NOR2_X1 U448 ( .A1(B[53]), .A2(A[53]), .ZN(n128) );
  NAND2_X1 U449 ( .A1(n28), .A2(n29), .ZN(net447659) );
  NAND2_X1 U450 ( .A1(n102), .A2(n99), .ZN(n108) );
  OR2_X1 U451 ( .A1(B[61]), .A2(A[61]), .ZN(n112) );
  NAND2_X1 U452 ( .A1(B[61]), .A2(A[61]), .ZN(net447636) );
  OR2_X1 U453 ( .A1(B[60]), .A2(A[60]), .ZN(n29) );
  NAND2_X1 U454 ( .A1(A[45]), .A2(B[45]), .ZN(n190) );
  OAI211_X1 U455 ( .C1(n200), .C2(n201), .A(n202), .B(n203), .ZN(n49) );
  AOI21_X1 U456 ( .B1(n256), .B2(n57), .A(n562), .ZN(n253) );
  NAND2_X1 U457 ( .A1(A[50]), .A2(B[50]), .ZN(n164) );
  INV_X1 U458 ( .A(n190), .ZN(n552) );
  XNOR2_X1 U459 ( .A(n518), .B(n314), .ZN(SUM[34]) );
  NAND2_X1 U460 ( .A1(n518), .A2(n304), .ZN(n312) );
  NAND2_X1 U461 ( .A1(n207), .A2(n239), .ZN(n240) );
  AND3_X1 U462 ( .A1(n220), .A2(n207), .A3(n208), .ZN(n202) );
  NAND2_X1 U463 ( .A1(n534), .A2(n177), .ZN(n172) );
  NAND2_X1 U464 ( .A1(B[56]), .A2(A[56]), .ZN(net447667) );
  AND2_X1 U465 ( .A1(net447669), .A2(n6), .ZN(net447695) );
  AND2_X1 U466 ( .A1(A[59]), .A2(B[59]), .ZN(net535350) );
  XNOR2_X1 U467 ( .A(n193), .B(n195), .ZN(SUM[49]) );
  NAND2_X1 U468 ( .A1(n272), .A2(n270), .ZN(n292) );
  NAND2_X1 U469 ( .A1(n2), .A2(n269), .ZN(n266) );
  NAND2_X1 U470 ( .A1(n272), .A2(n273), .ZN(n271) );
  NOR2_X1 U471 ( .A1(n531), .A2(n532), .ZN(n149) );
  AOI21_X1 U472 ( .B1(n121), .B2(n120), .A(n54), .ZN(n148) );
  OAI21_X1 U473 ( .B1(net447660), .B2(n522), .A(net447662), .ZN(net447656) );
  XNOR2_X1 U474 ( .A(n148), .B(n149), .ZN(SUM[53]) );
  XNOR2_X1 U475 ( .A(n109), .B(n111), .ZN(SUM[62]) );
  OAI21_X1 U476 ( .B1(n520), .B2(n541), .A(net447636), .ZN(n109) );
  XNOR2_X1 U477 ( .A(n519), .B(n260), .ZN(SUM[41]) );
  OAI21_X1 U478 ( .B1(n519), .B2(n61), .A(n250), .ZN(n40) );
  OAI21_X1 U479 ( .B1(n519), .B2(n61), .A(n250), .ZN(n256) );
  AOI21_X1 U480 ( .B1(n536), .B2(net447664), .A(net535350), .ZN(net447662) );
  NAND2_X1 U481 ( .A1(n153), .A2(n159), .ZN(n194) );
  NAND2_X1 U482 ( .A1(net447636), .A2(n112), .ZN(n113) );
  OAI211_X1 U483 ( .C1(net447666), .C2(net447667), .A(net447668), .B(net447669), .ZN(net447664) );
  NAND2_X1 U484 ( .A1(net447702), .A2(net447667), .ZN(net447701) );
  OAI21_X1 U485 ( .B1(net447666), .B2(net447667), .A(net447668), .ZN(net447692) );
  OAI211_X1 U486 ( .C1(n70), .C2(n223), .A(n214), .B(n215), .ZN(n275) );
  NAND2_X1 U487 ( .A1(n297), .A2(n298), .ZN(n214) );
  OAI211_X1 U488 ( .C1(n128), .C2(n129), .A(n130), .B(n131), .ZN(n127) );
  NAND2_X1 U489 ( .A1(n129), .A2(n146), .ZN(n145) );
  NAND2_X1 U490 ( .A1(net447673), .A2(net447674), .ZN(net447693) );
  NAND2_X1 U491 ( .A1(net447672), .A2(net447673), .ZN(net447702) );
  AOI21_X1 U492 ( .B1(n143), .B2(n502), .A(n145), .ZN(n141) );
  AOI21_X1 U493 ( .B1(n134), .B2(n60), .A(n531), .ZN(n137) );
  XNOR2_X1 U494 ( .A(n349), .B(n350), .ZN(SUM[30]) );
  NAND2_X1 U495 ( .A1(n349), .A2(n328), .ZN(n348) );
  INV_X1 U496 ( .A(net447676), .ZN(n537) );
  OAI211_X1 U497 ( .C1(A[45]), .C2(B[45]), .A(A[44]), .B(B[44]), .ZN(n189) );
  NAND2_X1 U498 ( .A1(B[44]), .A2(A[44]), .ZN(n239) );
  INV_X1 U499 ( .A(net447675), .ZN(n543) );
  NAND2_X1 U500 ( .A1(net447692), .A2(net447675), .ZN(net447691) );
  XNOR2_X1 U501 ( .A(net447672), .B(net447705), .ZN(SUM[56]) );
  AND2_X1 U502 ( .A1(A[55]), .A2(B[55]), .ZN(n74) );
  OR2_X1 U503 ( .A1(A[55]), .A2(B[55]), .ZN(n122) );
  NAND2_X1 U504 ( .A1(net447667), .A2(net447673), .ZN(net447705) );
  AOI21_X1 U505 ( .B1(n550), .B2(n220), .A(n552), .ZN(n232) );
  AOI21_X1 U506 ( .B1(n230), .B2(n208), .A(n73), .ZN(n228) );
  XNOR2_X1 U507 ( .A(n179), .B(n63), .ZN(SUM[50]) );
  XNOR2_X1 U508 ( .A(n289), .B(n65), .ZN(SUM[38]) );
  AOI21_X1 U509 ( .B1(n289), .B2(n224), .A(n547), .ZN(n285) );
  OAI21_X1 U510 ( .B1(n33), .B2(n557), .A(n272), .ZN(n289) );
  INV_X1 U511 ( .A(n106), .ZN(n538) );
  AOI21_X1 U512 ( .B1(n106), .B2(n109), .A(n539), .ZN(n107) );
  NAND2_X1 U513 ( .A1(n106), .A2(n103), .ZN(n111) );
  NAND2_X1 U514 ( .A1(B[63]), .A2(A[63]), .ZN(n102) );
  OAI211_X1 U515 ( .C1(n529), .C2(n163), .A(n171), .B(n164), .ZN(n144) );
  XNOR2_X1 U516 ( .A(net447701), .B(net447700), .ZN(SUM[57]) );
  INV_X1 U517 ( .A(n19), .ZN(n519) );
  NAND2_X1 U518 ( .A1(A[57]), .A2(B[57]), .ZN(net447668) );
  XNOR2_X1 U519 ( .A(n132), .B(n64), .ZN(SUM[55]) );
  AOI21_X1 U521 ( .B1(n134), .B2(n133), .A(n135), .ZN(n132) );
  AOI21_X1 U522 ( .B1(n530), .B2(n182), .A(n528), .ZN(n179) );
  OAI21_X1 U523 ( .B1(n506), .B2(B[47]), .A(n186), .ZN(n229) );
  NAND2_X1 U524 ( .A1(n506), .A2(B[47]), .ZN(n186) );
  INV_X1 U526 ( .A(A[47]), .ZN(n554) );
  OR2_X1 U528 ( .A1(A[47]), .A2(B[47]), .ZN(n32) );
  OR2_X1 U529 ( .A1(B[59]), .A2(A[59]), .ZN(net447676) );
  NAND4_X1 U530 ( .A1(n318), .A2(n319), .A3(n320), .A4(n321), .ZN(n305) );
  XNOR2_X1 U531 ( .A(n137), .B(n138), .ZN(SUM[54]) );
  AND2_X1 U532 ( .A1(A[52]), .A2(B[52]), .ZN(n54) );
  NAND2_X1 U534 ( .A1(A[52]), .A2(B[52]), .ZN(n129) );
  NOR2_X1 U535 ( .A1(n74), .A2(n498), .ZN(n64) );
  NOR2_X1 U536 ( .A1(n62), .A2(n68), .ZN(n126) );
  XNOR2_X1 U538 ( .A(n253), .B(n254), .ZN(SUM[43]) );
  OAI21_X1 U539 ( .B1(n263), .B2(n559), .A(n264), .ZN(n19) );
  NAND2_X1 U540 ( .A1(A[37]), .A2(B[37]), .ZN(n272) );
  AOI21_X1 U541 ( .B1(net447689), .B2(net537785), .A(net447690), .ZN(net447684) );
  NAND2_X1 U542 ( .A1(net447691), .A2(net447669), .ZN(net447690) );
  NOR2_X1 U543 ( .A1(net447693), .A2(n543), .ZN(net447689) );
  XNOR2_X1 U544 ( .A(net447684), .B(net447685), .ZN(SUM[59]) );
  NAND2_X1 U545 ( .A1(n194), .A2(n163), .ZN(n193) );
  INV_X1 U546 ( .A(n163), .ZN(n533) );
  NAND2_X1 U547 ( .A1(n163), .A2(n186), .ZN(n178) );
  XNOR2_X1 U548 ( .A(n507), .B(n240), .ZN(SUM[44]) );
  AOI21_X1 U550 ( .B1(n207), .B2(n507), .A(n550), .ZN(n237) );
  NAND2_X1 U551 ( .A1(n233), .A2(n232), .ZN(n230) );
  NAND2_X1 U552 ( .A1(n18), .A2(n118), .ZN(net447672) );
  NOR2_X1 U553 ( .A1(B[54]), .A2(A[54]), .ZN(n68) );
  NAND2_X1 U554 ( .A1(A[54]), .A2(B[54]), .ZN(n130) );
  AOI21_X1 U555 ( .B1(n127), .B2(n126), .A(n74), .ZN(n7) );
  AOI21_X1 U556 ( .B1(n126), .B2(n127), .A(n74), .ZN(n18) );
  NAND2_X1 U557 ( .A1(n169), .A2(n158), .ZN(n168) );
  INV_X1 U558 ( .A(n158), .ZN(n527) );
  AND2_X1 U559 ( .A1(n157), .A2(n158), .ZN(n143) );
  NAND2_X1 U560 ( .A1(n157), .A2(n158), .ZN(n156) );
  XNOR2_X1 U561 ( .A(net447694), .B(net447695), .ZN(SUM[58]) );
  AOI21_X1 U562 ( .B1(n514), .B2(net537785), .A(net447692), .ZN(net447694) );
  AND4_X1 U563 ( .A1(n177), .A2(n174), .A3(n175), .A4(n186), .ZN(n45) );
  NAND4_X1 U564 ( .A1(n49), .A2(n175), .A3(n177), .A4(n186), .ZN(n153) );
  NAND2_X1 U565 ( .A1(n171), .A2(n160), .ZN(n195) );
  NAND2_X1 U566 ( .A1(n159), .A2(n160), .ZN(n155) );
  INV_X1 U567 ( .A(n160), .ZN(n529) );
  NAND2_X1 U568 ( .A1(n160), .A2(n159), .ZN(n170) );
  INV_X1 U569 ( .A(n23), .ZN(n518) );
  AOI21_X1 U570 ( .B1(n315), .B2(n307), .A(n563), .ZN(n23) );
  NAND2_X1 U571 ( .A1(n497), .A2(B[31]), .ZN(n321) );
  OR2_X1 U572 ( .A1(A[31]), .A2(B[31]), .ZN(n329) );
  XNOR2_X1 U573 ( .A(n113), .B(net447653), .ZN(SUM[61]) );
  INV_X1 U574 ( .A(net447653), .ZN(n520) );
  INV_X1 U575 ( .A(n24), .ZN(n536) );
  NAND2_X1 U576 ( .A1(n141), .A2(n42), .ZN(n134) );
  NOR2_X1 U577 ( .A1(A[55]), .A2(B[55]), .ZN(n62) );
  INV_X1 U578 ( .A(net447656), .ZN(n521) );
  XNOR2_X1 U579 ( .A(net447659), .B(net447656), .ZN(SUM[60]) );
  OAI22_X1 U580 ( .A1(A[59]), .A2(B[59]), .B1(B[58]), .B2(A[58]), .ZN(n24) );
  OR2_X1 U581 ( .A1(A[58]), .A2(B[58]), .ZN(net447675) );
  OR2_X1 U582 ( .A1(B[58]), .A2(A[58]), .ZN(n6) );
  NAND2_X1 U583 ( .A1(A[58]), .A2(B[58]), .ZN(net447669) );
  NAND2_X1 U584 ( .A1(B[60]), .A2(A[60]), .ZN(n28) );
endmodule


module RCA_NBIT64_4 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_4_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_3_DW01_add_5 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net446593, net446587, net446564, net446543, net446539, net446536,
         net446535, net446534, net446530, net446526, net446521, net446520,
         net446519, net446511, net446502, net446501, net446484, net535419,
         net537284, net538437, net538658, net446508, net446490, net446522,
         net537208, net446594, net446517, net446516, net446514, net446513,
         net446512, net446509, net446505, net446491, n1, n2, n4, n6, n8, n9,
         n10, n14, n16, n17, n18, n20, n21, n23, n25, n27, n28, n30, n31, n35,
         n36, n37, n38, n41, n42, n45, n50, n51, n52, n54, n56, n57, n59, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n107,
         n108, n109, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n135, n137, n138, n140, n141, n144, n145, n146,
         n148, n149, n150, n152, n153, n154, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n174,
         n175, n177, n178, n179, n180, n181, n182, n183, n184, n185, n188,
         n189, n191, n192, n193, n195, n196, n197, n198, n200, n202, n203,
         n206, n207, n208, n211, n212, n213, n214, n215, n216, n217, n219,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n234,
         n237, n239, n240, n241, n242, n243, n244, n245, n246, n248, n249,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n272, n274, n276,
         n277, n278, n279, n280, n281, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n321, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n347, n348, n349,
         n350, n352, n354, n355, n356, n359, n360, n361, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n375, n376, n377, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n396, n397, n399, n400, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n421, n423, n424, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n448, n449, n450, n451, n452, n453, n454,
         n455, n457, n459, n460, n461, n462, n463, n466, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n502, n503, n504, n505, n508,
         n509, n510, n511, n512, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608;

  NAND3_X1 U40 ( .A1(n254), .A2(n203), .A3(n253), .ZN(n25) );
  OR2_X2 U48 ( .A1(B[44]), .A2(A[44]), .ZN(n234) );
  OR2_X2 U49 ( .A1(A[42]), .A2(B[42]), .ZN(n263) );
  OR2_X2 U123 ( .A1(A[58]), .A2(B[58]), .ZN(net446520) );
  OR2_X2 U359 ( .A1(B[45]), .A2(A[45]), .ZN(n202) );
  NAND3_X1 U522 ( .A1(n121), .A2(n120), .A3(n131), .ZN(n103) );
  NAND3_X1 U523 ( .A1(n524), .A2(B[52]), .A3(n516), .ZN(n120) );
  NAND3_X1 U528 ( .A1(A[49]), .A2(B[48]), .A3(A[48]), .ZN(n162) );
  NAND3_X1 U529 ( .A1(B[49]), .A2(A[48]), .A3(B[48]), .ZN(n161) );
  NAND3_X1 U531 ( .A1(n177), .A2(n200), .A3(n178), .ZN(n171) );
  NAND3_X1 U532 ( .A1(n183), .A2(n184), .A3(n185), .ZN(n182) );
  NAND3_X1 U543 ( .A1(n206), .A2(n207), .A3(n208), .ZN(n179) );
  NAND3_X1 U544 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n207) );
  NAND3_X1 U551 ( .A1(n237), .A2(n542), .A3(n239), .ZN(n225) );
  NAND3_X1 U553 ( .A1(n245), .A2(n202), .A3(n230), .ZN(n244) );
  NAND3_X1 U558 ( .A1(n254), .A2(n203), .A3(n253), .ZN(n245) );
  NAND3_X1 U560 ( .A1(n215), .A2(n216), .A3(n212), .ZN(n257) );
  NAND3_X1 U561 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n212) );
  NAND3_X1 U562 ( .A1(n9), .A2(n267), .A3(n266), .ZN(n255) );
  NAND3_X1 U574 ( .A1(n287), .A2(n288), .A3(n237), .ZN(n286) );
  NAND3_X1 U575 ( .A1(n239), .A2(n45), .A3(n294), .ZN(n278) );
  NAND3_X1 U612 ( .A1(n490), .A2(n491), .A3(n492), .ZN(n489) );
  NAND3_X1 U613 ( .A1(n493), .A2(n65), .A3(n494), .ZN(n490) );
  NAND3_X1 U618 ( .A1(n504), .A2(n75), .A3(n74), .ZN(n503) );
  NAND3_X1 U619 ( .A1(n83), .A2(n505), .A3(n78), .ZN(n504) );
  OR2_X2 U89 ( .A1(B[60]), .A2(A[60]), .ZN(net446505) );
  OR2_X2 U130 ( .A1(B[48]), .A2(A[48]), .ZN(n166) );
  INV_X1 U2 ( .A(n562), .ZN(n515) );
  OR2_X1 U3 ( .A1(A[43]), .A2(B[43]), .ZN(n256) );
  OR2_X1 U4 ( .A1(A[41]), .A2(B[41]), .ZN(n261) );
  AND2_X1 U5 ( .A1(n508), .A2(n441), .ZN(SUM[0]) );
  INV_X1 U6 ( .A(n526), .ZN(net446491) );
  OR2_X2 U7 ( .A1(A[49]), .A2(B[49]), .ZN(n167) );
  CLKBUF_X1 U8 ( .A(A[52]), .Z(n516) );
  AND2_X1 U9 ( .A1(n256), .A2(n234), .ZN(n517) );
  NAND2_X1 U10 ( .A1(n159), .A2(n160), .ZN(n518) );
  CLKBUF_X1 U11 ( .A(n41), .Z(n519) );
  AND2_X1 U12 ( .A1(A[60]), .A2(B[60]), .ZN(n526) );
  INV_X1 U13 ( .A(n121), .ZN(n574) );
  INV_X1 U14 ( .A(n545), .ZN(n520) );
  NAND2_X1 U15 ( .A1(n257), .A2(n517), .ZN(n253) );
  OR2_X2 U16 ( .A1(B[38]), .A2(A[38]), .ZN(n237) );
  AND2_X1 U17 ( .A1(n521), .A2(n234), .ZN(n228) );
  NOR3_X1 U18 ( .A1(n532), .A2(n225), .A3(n533), .ZN(n521) );
  OR2_X1 U19 ( .A1(A[54]), .A2(B[54]), .ZN(n133) );
  NAND3_X1 U20 ( .A1(n206), .A2(n207), .A3(n208), .ZN(n522) );
  INV_X1 U21 ( .A(n524), .ZN(n523) );
  OR2_X1 U22 ( .A1(A[53]), .A2(B[53]), .ZN(n524) );
  OR2_X1 U23 ( .A1(A[50]), .A2(B[50]), .ZN(n1) );
  AND4_X2 U24 ( .A1(n177), .A2(n180), .A3(n179), .A4(n200), .ZN(n52) );
  AND2_X1 U25 ( .A1(n14), .A2(n140), .ZN(n525) );
  AND2_X1 U26 ( .A1(n127), .A2(n525), .ZN(n62) );
  OR2_X1 U27 ( .A1(B[55]), .A2(A[55]), .ZN(n10) );
  OR2_X2 U28 ( .A1(A[61]), .A2(B[61]), .ZN(net538437) );
  XNOR2_X1 U29 ( .A(n529), .B(n527), .ZN(SUM[56]) );
  NAND2_X1 U30 ( .A1(n51), .A2(net446534), .ZN(n527) );
  XOR2_X1 U31 ( .A(n52), .B(n528), .Z(SUM[48]) );
  NAND2_X1 U32 ( .A1(n166), .A2(n198), .ZN(n528) );
  INV_X1 U33 ( .A(n399), .ZN(n584) );
  INV_X1 U34 ( .A(n439), .ZN(n593) );
  AOI21_X1 U35 ( .B1(n99), .B2(net446511), .A(net446530), .ZN(net538658) );
  NOR2_X1 U36 ( .A1(n224), .A2(n225), .ZN(n217) );
  INV_X1 U37 ( .A(n223), .ZN(n541) );
  NOR3_X1 U38 ( .A1(n547), .A2(n549), .A3(n543), .ZN(n219) );
  NOR2_X1 U39 ( .A1(n543), .A2(n549), .ZN(n266) );
  NAND2_X1 U41 ( .A1(n278), .A2(n223), .ZN(n267) );
  NOR2_X1 U42 ( .A1(n547), .A2(n545), .ZN(n232) );
  OAI21_X1 U43 ( .B1(n606), .B2(n475), .A(n472), .ZN(n68) );
  OAI21_X1 U44 ( .B1(n593), .B2(n361), .A(n589), .ZN(n413) );
  INV_X1 U45 ( .A(n352), .ZN(n589) );
  OAI21_X1 U46 ( .B1(n588), .B2(n355), .A(n354), .ZN(n399) );
  INV_X1 U47 ( .A(n413), .ZN(n588) );
  AOI21_X1 U50 ( .B1(n471), .B2(n472), .A(n473), .ZN(n466) );
  NAND2_X1 U51 ( .A1(n601), .A2(n474), .ZN(n471) );
  INV_X1 U52 ( .A(n475), .ZN(n601) );
  NAND2_X1 U53 ( .A1(n452), .A2(n453), .ZN(n439) );
  OAI21_X1 U54 ( .B1(n466), .B2(n598), .A(n16), .ZN(n452) );
  AOI21_X1 U55 ( .B1(n454), .B2(n455), .A(n594), .ZN(n453) );
  INV_X1 U56 ( .A(n470), .ZN(n598) );
  NAND4_X1 U57 ( .A1(n59), .A2(n590), .A3(n579), .A4(n356), .ZN(n335) );
  INV_X1 U58 ( .A(n361), .ZN(n590) );
  INV_X1 U59 ( .A(n350), .ZN(n579) );
  NOR2_X1 U60 ( .A1(n593), .A2(n355), .ZN(n356) );
  NAND2_X1 U61 ( .A1(n487), .A2(n470), .ZN(n485) );
  NAND2_X1 U62 ( .A1(n597), .A2(n68), .ZN(n487) );
  INV_X1 U63 ( .A(n473), .ZN(n597) );
  INV_X1 U64 ( .A(n474), .ZN(n606) );
  INV_X1 U65 ( .A(n355), .ZN(n583) );
  NOR2_X1 U66 ( .A1(n85), .A2(n567), .ZN(SUM[64]) );
  INV_X1 U67 ( .A(n354), .ZN(n585) );
  NAND2_X1 U68 ( .A1(n153), .A2(n152), .ZN(n158) );
  NAND2_X1 U69 ( .A1(n237), .A2(n292), .ZN(n309) );
  NAND3_X1 U70 ( .A1(n102), .A2(net446539), .A3(n112), .ZN(n529) );
  NOR2_X1 U71 ( .A1(net446594), .A2(net446539), .ZN(net446593) );
  NAND2_X1 U72 ( .A1(n317), .A2(n324), .ZN(n330) );
  NAND2_X1 U73 ( .A1(n263), .A2(n216), .ZN(n274) );
  NAND2_X1 U74 ( .A1(n202), .A2(n183), .ZN(n252) );
  XNOR2_X1 U75 ( .A(n196), .B(n197), .ZN(SUM[49]) );
  NOR2_X1 U76 ( .A1(n557), .A2(n558), .ZN(n197) );
  AOI21_X1 U77 ( .B1(n168), .B2(n166), .A(n556), .ZN(n196) );
  NOR2_X1 U78 ( .A1(n573), .A2(n572), .ZN(n150) );
  INV_X1 U79 ( .A(n131), .ZN(n573) );
  AOI21_X1 U80 ( .B1(n171), .B2(n170), .A(n172), .ZN(n169) );
  AND3_X1 U81 ( .A1(n167), .A2(n1), .A3(n166), .ZN(n170) );
  NAND2_X1 U82 ( .A1(n180), .A2(n6), .ZN(n241) );
  NAND2_X1 U83 ( .A1(n244), .A2(n243), .ZN(n242) );
  XNOR2_X1 U84 ( .A(n109), .B(net537284), .ZN(SUM[59]) );
  INV_X1 U85 ( .A(net446535), .ZN(n571) );
  XOR2_X1 U86 ( .A(n530), .B(n368), .Z(SUM[29]) );
  NAND2_X1 U87 ( .A1(n345), .A2(n360), .ZN(n530) );
  AND3_X1 U88 ( .A1(n232), .A2(n202), .A3(n211), .ZN(n231) );
  OAI211_X1 U90 ( .C1(n560), .C2(n101), .A(n102), .B(net446539), .ZN(net446511) );
  INV_X1 U91 ( .A(n103), .ZN(n560) );
  OAI21_X1 U92 ( .B1(n549), .B2(n278), .A(n279), .ZN(n276) );
  INV_X1 U93 ( .A(n265), .ZN(n548) );
  AND2_X1 U94 ( .A1(n283), .A2(n239), .ZN(n280) );
  OAI211_X1 U95 ( .C1(n538), .C2(n323), .A(n324), .B(n325), .ZN(n318) );
  NOR2_X1 U96 ( .A1(n544), .A2(n545), .ZN(n270) );
  AOI21_X1 U97 ( .B1(n272), .B2(n263), .A(n546), .ZN(n269) );
  INV_X1 U98 ( .A(n215), .ZN(n544) );
  AND2_X1 U99 ( .A1(net446539), .A2(n10), .ZN(n57) );
  NAND2_X1 U100 ( .A1(n146), .A2(n131), .ZN(n145) );
  XNOR2_X1 U101 ( .A(n248), .B(n249), .ZN(SUM[46]) );
  NOR2_X1 U102 ( .A1(n552), .A2(n554), .ZN(n249) );
  AOI21_X1 U103 ( .B1(n202), .B2(n245), .A(n551), .ZN(n248) );
  INV_X1 U104 ( .A(n183), .ZN(n551) );
  XOR2_X1 U105 ( .A(n154), .B(n531), .Z(SUM[53]) );
  OR2_X1 U106 ( .A1(n574), .A2(n523), .ZN(n531) );
  NAND2_X1 U107 ( .A1(n558), .A2(n1), .ZN(n175) );
  OAI21_X1 U108 ( .B1(n536), .B2(n368), .A(n345), .ZN(n366) );
  XNOR2_X1 U109 ( .A(n188), .B(n189), .ZN(SUM[50]) );
  NOR2_X1 U110 ( .A1(n576), .A2(n575), .ZN(n189) );
  AOI21_X1 U111 ( .B1(n191), .B2(n168), .A(n192), .ZN(n188) );
  AOI21_X1 U112 ( .B1(n539), .B2(n318), .A(n540), .ZN(n224) );
  INV_X1 U113 ( .A(n321), .ZN(n540) );
  INV_X1 U114 ( .A(n31), .ZN(n539) );
  XNOR2_X1 U115 ( .A(n334), .B(n28), .ZN(SUM[32]) );
  NAND2_X1 U116 ( .A1(n315), .A2(n323), .ZN(n334) );
  INV_X1 U117 ( .A(n240), .ZN(n542) );
  OAI21_X1 U118 ( .B1(n535), .B2(n543), .A(n264), .ZN(n272) );
  INV_X1 U119 ( .A(n276), .ZN(n535) );
  XNOR2_X1 U120 ( .A(n326), .B(n327), .ZN(SUM[35]) );
  NAND2_X1 U121 ( .A1(n328), .A2(n324), .ZN(n326) );
  XNOR2_X1 U122 ( .A(n364), .B(n363), .ZN(SUM[31]) );
  NAND2_X1 U124 ( .A1(n343), .A2(n338), .ZN(n363) );
  NAND2_X1 U125 ( .A1(n365), .A2(n344), .ZN(n364) );
  NAND2_X1 U126 ( .A1(n366), .A2(n342), .ZN(n365) );
  XNOR2_X1 U127 ( .A(n313), .B(n45), .ZN(SUM[36]) );
  NAND2_X1 U128 ( .A1(n296), .A2(n290), .ZN(n313) );
  NOR2_X1 U129 ( .A1(n578), .A2(n240), .ZN(n294) );
  INV_X1 U131 ( .A(n237), .ZN(n578) );
  XNOR2_X1 U132 ( .A(n276), .B(n277), .ZN(SUM[41]) );
  NAND2_X1 U133 ( .A1(n264), .A2(n261), .ZN(n277) );
  XNOR2_X1 U134 ( .A(n284), .B(n267), .ZN(SUM[40]) );
  NAND2_X1 U135 ( .A1(n283), .A2(n265), .ZN(n284) );
  XNOR2_X1 U136 ( .A(n258), .B(n259), .ZN(SUM[44]) );
  NAND2_X1 U137 ( .A1(n234), .A2(n203), .ZN(n258) );
  NAND2_X1 U138 ( .A1(n255), .A2(n260), .ZN(n259) );
  XNOR2_X1 U139 ( .A(n23), .B(n311), .ZN(SUM[37]) );
  NAND2_X1 U140 ( .A1(n287), .A2(n289), .ZN(n311) );
  NAND2_X1 U141 ( .A1(n312), .A2(n290), .ZN(n23) );
  XNOR2_X1 U142 ( .A(n377), .B(n376), .ZN(SUM[28]) );
  NAND2_X1 U143 ( .A1(n359), .A2(n347), .ZN(n377) );
  XNOR2_X1 U144 ( .A(n332), .B(n331), .ZN(SUM[33]) );
  NAND2_X1 U145 ( .A1(n316), .A2(n325), .ZN(n332) );
  NAND2_X1 U146 ( .A1(n333), .A2(n323), .ZN(n331) );
  XNOR2_X1 U147 ( .A(n366), .B(n367), .ZN(SUM[30]) );
  NAND2_X1 U148 ( .A1(n342), .A2(n344), .ZN(n367) );
  XNOR2_X1 U149 ( .A(n389), .B(n390), .ZN(SUM[27]) );
  NAND2_X1 U150 ( .A1(n382), .A2(n391), .ZN(n389) );
  NAND2_X1 U151 ( .A1(n380), .A2(n381), .ZN(n390) );
  NAND2_X1 U152 ( .A1(n392), .A2(n385), .ZN(n391) );
  XNOR2_X1 U153 ( .A(n397), .B(n396), .ZN(SUM[25]) );
  NAND2_X1 U154 ( .A1(n383), .A2(n386), .ZN(n397) );
  XNOR2_X1 U155 ( .A(n393), .B(n392), .ZN(SUM[26]) );
  NAND2_X1 U156 ( .A1(n385), .A2(n382), .ZN(n393) );
  NAND4_X1 U157 ( .A1(n177), .A2(n522), .A3(n200), .A4(n180), .ZN(n168) );
  NOR2_X1 U158 ( .A1(n226), .A2(n227), .ZN(n206) );
  INV_X1 U159 ( .A(net446534), .ZN(n566) );
  OAI21_X1 U160 ( .B1(n21), .B2(n538), .A(n325), .ZN(n329) );
  AND2_X1 U161 ( .A1(n333), .A2(n323), .ZN(n21) );
  NOR2_X1 U162 ( .A1(n104), .A2(net446543), .ZN(n99) );
  NAND2_X1 U163 ( .A1(net446522), .A2(n565), .ZN(net446543) );
  XNOR2_X1 U164 ( .A(n306), .B(n305), .ZN(SUM[39]) );
  NAND2_X1 U165 ( .A1(n291), .A2(n239), .ZN(n305) );
  NAND2_X1 U166 ( .A1(n307), .A2(n292), .ZN(n306) );
  INV_X1 U167 ( .A(n261), .ZN(n543) );
  OAI21_X1 U168 ( .B1(n339), .B2(n340), .A(n341), .ZN(n337) );
  NOR2_X1 U169 ( .A1(n536), .A2(n347), .ZN(n339) );
  NAND2_X1 U170 ( .A1(n344), .A2(n345), .ZN(n340) );
  AND2_X1 U171 ( .A1(n343), .A2(n342), .ZN(n341) );
  INV_X1 U172 ( .A(n283), .ZN(n549) );
  AND2_X1 U173 ( .A1(n291), .A2(n292), .ZN(n285) );
  NAND2_X1 U174 ( .A1(n289), .A2(n290), .ZN(n288) );
  AND2_X1 U175 ( .A1(n522), .A2(n180), .ZN(n178) );
  OAI21_X1 U176 ( .B1(n584), .B2(n350), .A(n20), .ZN(n376) );
  OAI21_X1 U177 ( .B1(n17), .B2(n379), .A(n380), .ZN(n20) );
  NAND2_X1 U178 ( .A1(n264), .A2(n265), .ZN(n262) );
  NOR2_X1 U179 ( .A1(n246), .A2(n554), .ZN(n243) );
  NOR2_X1 U180 ( .A1(n552), .A2(n183), .ZN(n246) );
  NAND3_X1 U181 ( .A1(n519), .A2(n317), .A3(n54), .ZN(n532) );
  OR2_X1 U182 ( .A1(n543), .A2(n549), .ZN(n533) );
  NOR2_X1 U183 ( .A1(n555), .A2(n557), .ZN(n191) );
  INV_X1 U184 ( .A(n166), .ZN(n555) );
  XNOR2_X1 U185 ( .A(n419), .B(n421), .ZN(SUM[21]) );
  NOR2_X1 U186 ( .A1(n587), .A2(n586), .ZN(n421) );
  INV_X1 U187 ( .A(n410), .ZN(n587) );
  AND2_X1 U188 ( .A1(n375), .A2(n347), .ZN(n368) );
  NAND2_X1 U189 ( .A1(n376), .A2(n359), .ZN(n375) );
  NAND2_X1 U190 ( .A1(n239), .A2(n281), .ZN(n223) );
  NAND2_X1 U191 ( .A1(n381), .A2(n382), .ZN(n379) );
  NAND2_X1 U192 ( .A1(n181), .A2(n182), .ZN(n200) );
  AND2_X1 U193 ( .A1(n6), .A2(n8), .ZN(n181) );
  NAND2_X1 U194 ( .A1(n605), .A2(n553), .ZN(n8) );
  NAND2_X1 U195 ( .A1(n296), .A2(n287), .ZN(n240) );
  NAND2_X1 U196 ( .A1(n293), .A2(n296), .ZN(n312) );
  INV_X1 U197 ( .A(n318), .ZN(n537) );
  AOI21_X1 U198 ( .B1(n310), .B2(n287), .A(n577), .ZN(n30) );
  INV_X1 U199 ( .A(n289), .ZN(n577) );
  NAND2_X1 U200 ( .A1(n312), .A2(n290), .ZN(n310) );
  INV_X1 U201 ( .A(n193), .ZN(n558) );
  NAND2_X1 U202 ( .A1(n556), .A2(n167), .ZN(n174) );
  NAND2_X1 U203 ( .A1(n229), .A2(n315), .ZN(n333) );
  INV_X1 U204 ( .A(n167), .ZN(n557) );
  NAND2_X1 U205 ( .A1(n135), .A2(n10), .ZN(n125) );
  INV_X1 U206 ( .A(net446594), .ZN(n565) );
  INV_X1 U207 ( .A(n185), .ZN(n554) );
  INV_X1 U208 ( .A(n263), .ZN(n547) );
  INV_X1 U209 ( .A(n408), .ZN(n586) );
  AND4_X1 U210 ( .A1(n343), .A2(n360), .A3(n342), .A4(n359), .ZN(n59) );
  NAND2_X1 U211 ( .A1(n174), .A2(n193), .ZN(n192) );
  INV_X1 U212 ( .A(n360), .ZN(n536) );
  INV_X1 U213 ( .A(n316), .ZN(n538) );
  INV_X1 U214 ( .A(n198), .ZN(n556) );
  AND3_X1 U215 ( .A1(n120), .A2(n121), .A3(n131), .ZN(n61) );
  NAND2_X1 U216 ( .A1(n42), .A2(n234), .ZN(n254) );
  AND3_X1 U217 ( .A1(n268), .A2(n267), .A3(n266), .ZN(n42) );
  INV_X1 U218 ( .A(net446505), .ZN(n569) );
  NAND2_X1 U219 ( .A1(n59), .A2(n348), .ZN(n336) );
  OAI21_X1 U220 ( .B1(n349), .B2(n350), .A(n2), .ZN(n348) );
  AOI21_X1 U221 ( .B1(n583), .B2(n352), .A(n585), .ZN(n349) );
  OAI21_X1 U222 ( .B1(n17), .B2(n379), .A(n380), .ZN(n2) );
  INV_X1 U223 ( .A(n1), .ZN(n575) );
  NAND2_X1 U224 ( .A1(n550), .A2(n202), .ZN(n184) );
  INV_X1 U225 ( .A(n203), .ZN(n550) );
  INV_X1 U226 ( .A(n216), .ZN(n546) );
  AND2_X1 U227 ( .A1(n153), .A2(n524), .ZN(n14) );
  AND2_X1 U228 ( .A1(n316), .A2(n315), .ZN(n54) );
  NAND2_X1 U229 ( .A1(n56), .A2(net535419), .ZN(n111) );
  AND2_X1 U230 ( .A1(n102), .A2(n112), .ZN(n56) );
  INV_X1 U231 ( .A(n152), .ZN(n559) );
  AND2_X1 U232 ( .A1(n215), .A2(n216), .ZN(n214) );
  XNOR2_X1 U233 ( .A(n442), .B(n443), .ZN(SUM[19]) );
  NAND2_X1 U234 ( .A1(n433), .A2(n444), .ZN(n442) );
  NAND2_X1 U235 ( .A1(n428), .A2(n430), .ZN(n443) );
  NAND2_X1 U236 ( .A1(n445), .A2(n429), .ZN(n444) );
  XNOR2_X1 U237 ( .A(n476), .B(n477), .ZN(SUM[15]) );
  NAND2_X1 U238 ( .A1(n478), .A2(n461), .ZN(n477) );
  NAND2_X1 U239 ( .A1(n457), .A2(n463), .ZN(n476) );
  NAND2_X1 U240 ( .A1(n462), .A2(n479), .ZN(n478) );
  XNOR2_X1 U241 ( .A(n414), .B(n415), .ZN(SUM[23]) );
  NAND2_X1 U242 ( .A1(n406), .A2(n416), .ZN(n415) );
  NAND2_X1 U243 ( .A1(n405), .A2(n404), .ZN(n414) );
  NAND2_X1 U244 ( .A1(n409), .A2(n417), .ZN(n416) );
  XNOR2_X1 U245 ( .A(n424), .B(n413), .ZN(SUM[20]) );
  NAND2_X1 U246 ( .A1(n412), .A2(n411), .ZN(n424) );
  XNOR2_X1 U247 ( .A(n400), .B(n399), .ZN(SUM[24]) );
  NAND2_X1 U248 ( .A1(n388), .A2(n387), .ZN(n400) );
  XNOR2_X1 U249 ( .A(n480), .B(n479), .ZN(SUM[14]) );
  NAND2_X1 U250 ( .A1(n462), .A2(n461), .ZN(n480) );
  XNOR2_X1 U251 ( .A(n418), .B(n417), .ZN(SUM[22]) );
  NAND2_X1 U252 ( .A1(n409), .A2(n406), .ZN(n418) );
  XNOR2_X1 U253 ( .A(n451), .B(n439), .ZN(SUM[16]) );
  NAND2_X1 U254 ( .A1(n436), .A2(n437), .ZN(n451) );
  XNOR2_X1 U255 ( .A(n446), .B(n445), .ZN(SUM[18]) );
  NAND2_X1 U256 ( .A1(n429), .A2(n433), .ZN(n446) );
  XNOR2_X1 U257 ( .A(n449), .B(n448), .ZN(SUM[17]) );
  NAND2_X1 U258 ( .A1(n438), .A2(n434), .ZN(n449) );
  XNOR2_X1 U259 ( .A(n483), .B(n482), .ZN(SUM[13]) );
  NAND2_X1 U260 ( .A1(n469), .A2(n460), .ZN(n483) );
  XNOR2_X1 U261 ( .A(n71), .B(n72), .ZN(SUM[7]) );
  NAND2_X1 U262 ( .A1(n75), .A2(n76), .ZN(n71) );
  NAND2_X1 U263 ( .A1(n73), .A2(n74), .ZN(n72) );
  NAND2_X1 U264 ( .A1(n77), .A2(n78), .ZN(n76) );
  XNOR2_X1 U265 ( .A(n297), .B(n298), .ZN(SUM[3]) );
  NAND2_X1 U266 ( .A1(n301), .A2(n302), .ZN(n297) );
  NAND2_X1 U267 ( .A1(n299), .A2(n300), .ZN(n298) );
  NAND2_X1 U268 ( .A1(n303), .A2(n304), .ZN(n302) );
  XNOR2_X1 U269 ( .A(n495), .B(n496), .ZN(SUM[11]) );
  NAND2_X1 U270 ( .A1(n491), .A2(n497), .ZN(n496) );
  NAND2_X1 U271 ( .A1(n492), .A2(n488), .ZN(n495) );
  NAND2_X1 U272 ( .A1(n494), .A2(n498), .ZN(n497) );
  XNOR2_X1 U273 ( .A(n440), .B(n608), .ZN(SUM[1]) );
  NAND2_X1 U274 ( .A1(n372), .A2(n371), .ZN(n440) );
  XNOR2_X1 U275 ( .A(n486), .B(n485), .ZN(SUM[12]) );
  NAND2_X1 U276 ( .A1(n468), .A2(n459), .ZN(n486) );
  XNOR2_X1 U277 ( .A(n67), .B(n68), .ZN(SUM[8]) );
  NAND2_X1 U278 ( .A1(n69), .A2(n70), .ZN(n67) );
  XNOR2_X1 U279 ( .A(n105), .B(n84), .ZN(SUM[5]) );
  NAND2_X1 U280 ( .A1(n83), .A2(n82), .ZN(n105) );
  XNOR2_X1 U281 ( .A(n63), .B(n64), .ZN(SUM[9]) );
  NAND2_X1 U282 ( .A1(n65), .A2(n66), .ZN(n63) );
  XNOR2_X1 U283 ( .A(n79), .B(n77), .ZN(SUM[6]) );
  NAND2_X1 U284 ( .A1(n78), .A2(n75), .ZN(n79) );
  XNOR2_X1 U285 ( .A(n499), .B(n498), .ZN(SUM[10]) );
  NAND2_X1 U286 ( .A1(n494), .A2(n491), .ZN(n499) );
  XNOR2_X1 U287 ( .A(n369), .B(n303), .ZN(SUM[2]) );
  NAND2_X1 U288 ( .A1(n304), .A2(n301), .ZN(n369) );
  XNOR2_X1 U289 ( .A(n195), .B(n474), .ZN(SUM[4]) );
  NAND2_X1 U290 ( .A1(n108), .A2(n107), .ZN(n195) );
  OAI21_X1 U291 ( .B1(n509), .B2(n510), .A(n300), .ZN(n474) );
  NAND2_X1 U292 ( .A1(n304), .A2(n299), .ZN(n510) );
  NOR2_X1 U293 ( .A1(n511), .A2(n512), .ZN(n509) );
  NAND2_X1 U294 ( .A1(n301), .A2(n371), .ZN(n512) );
  OAI21_X1 U295 ( .B1(n600), .B2(n599), .A(n66), .ZN(n498) );
  INV_X1 U296 ( .A(n64), .ZN(n600) );
  INV_X1 U297 ( .A(n65), .ZN(n599) );
  OAI21_X1 U298 ( .B1(n596), .B2(n595), .A(n460), .ZN(n479) );
  INV_X1 U299 ( .A(n482), .ZN(n596) );
  OAI21_X1 U300 ( .B1(n419), .B2(n586), .A(n410), .ZN(n417) );
  OAI21_X1 U301 ( .B1(n582), .B2(n584), .A(n387), .ZN(n396) );
  INV_X1 U302 ( .A(n388), .ZN(n582) );
  OAI21_X1 U303 ( .B1(n604), .B2(n606), .A(n107), .ZN(n84) );
  INV_X1 U304 ( .A(n108), .ZN(n604) );
  OAI21_X1 U305 ( .B1(n603), .B2(n602), .A(n82), .ZN(n77) );
  INV_X1 U306 ( .A(n83), .ZN(n602) );
  INV_X1 U307 ( .A(n84), .ZN(n603) );
  OAI21_X1 U308 ( .B1(n581), .B2(n580), .A(n386), .ZN(n392) );
  INV_X1 U309 ( .A(n383), .ZN(n580) );
  INV_X1 U310 ( .A(n396), .ZN(n581) );
  OAI21_X1 U311 ( .B1(n592), .B2(n591), .A(n434), .ZN(n445) );
  INV_X1 U312 ( .A(n448), .ZN(n592) );
  NAND4_X1 U313 ( .A1(n412), .A2(n408), .A3(n409), .A4(n404), .ZN(n355) );
  NAND4_X1 U314 ( .A1(n388), .A2(n383), .A3(n385), .A4(n380), .ZN(n350) );
  OAI21_X1 U315 ( .B1(n426), .B2(n427), .A(n428), .ZN(n352) );
  NAND2_X1 U316 ( .A1(n429), .A2(n430), .ZN(n427) );
  NOR2_X1 U317 ( .A1(n431), .A2(n432), .ZN(n426) );
  NAND2_X1 U318 ( .A1(n433), .A2(n434), .ZN(n432) );
  OAI21_X1 U319 ( .B1(n402), .B2(n403), .A(n404), .ZN(n354) );
  NAND2_X1 U320 ( .A1(n405), .A2(n406), .ZN(n403) );
  NOR2_X1 U321 ( .A1(n18), .A2(n407), .ZN(n402) );
  AND2_X1 U322 ( .A1(n410), .A2(n411), .ZN(n18) );
  NAND4_X1 U323 ( .A1(n437), .A2(n438), .A3(n429), .A4(n430), .ZN(n361) );
  NAND4_X1 U324 ( .A1(n108), .A2(n83), .A3(n78), .A4(n73), .ZN(n475) );
  NAND4_X1 U325 ( .A1(n65), .A2(n69), .A3(n494), .A4(n488), .ZN(n473) );
  OAI211_X1 U326 ( .C1(n595), .C2(n459), .A(n460), .B(n461), .ZN(n455) );
  AOI21_X1 U327 ( .B1(n88), .B2(net446484), .A(n89), .ZN(n85) );
  NOR2_X1 U328 ( .A1(n591), .A2(n436), .ZN(n431) );
  NOR2_X1 U329 ( .A1(n607), .A2(n441), .ZN(n511) );
  INV_X1 U330 ( .A(n372), .ZN(n607) );
  NAND2_X1 U331 ( .A1(n502), .A2(n70), .ZN(n64) );
  NAND2_X1 U332 ( .A1(n68), .A2(n69), .ZN(n502) );
  NAND2_X1 U333 ( .A1(n484), .A2(n459), .ZN(n482) );
  NAND2_X1 U334 ( .A1(n485), .A2(n468), .ZN(n484) );
  NAND2_X1 U335 ( .A1(n450), .A2(n436), .ZN(n448) );
  NAND2_X1 U336 ( .A1(n439), .A2(n437), .ZN(n450) );
  NAND2_X1 U337 ( .A1(n370), .A2(n371), .ZN(n303) );
  NAND2_X1 U338 ( .A1(n372), .A2(n608), .ZN(n370) );
  NAND2_X1 U339 ( .A1(n488), .A2(n489), .ZN(n470) );
  NAND2_X1 U340 ( .A1(n66), .A2(n70), .ZN(n493) );
  NAND2_X1 U341 ( .A1(n73), .A2(n503), .ZN(n472) );
  NAND2_X1 U342 ( .A1(n82), .A2(n107), .ZN(n505) );
  AND3_X1 U343 ( .A1(n383), .A2(n384), .A3(n385), .ZN(n17) );
  NAND2_X1 U344 ( .A1(n386), .A2(n387), .ZN(n384) );
  INV_X1 U345 ( .A(n441), .ZN(n608) );
  AND2_X1 U346 ( .A1(n423), .A2(n411), .ZN(n419) );
  NAND2_X1 U347 ( .A1(n413), .A2(n412), .ZN(n423) );
  INV_X1 U348 ( .A(n438), .ZN(n591) );
  INV_X1 U349 ( .A(n469), .ZN(n595) );
  NAND2_X1 U350 ( .A1(n408), .A2(n409), .ZN(n407) );
  AND4_X1 U351 ( .A1(n468), .A2(n469), .A3(n462), .A4(n463), .ZN(n16) );
  AND2_X1 U352 ( .A1(n463), .A2(n462), .ZN(n454) );
  INV_X1 U353 ( .A(n87), .ZN(n567) );
  INV_X1 U354 ( .A(n457), .ZN(n594) );
  NOR2_X1 U355 ( .A1(n516), .A2(B[52]), .ZN(n137) );
  NAND2_X1 U356 ( .A1(A[55]), .A2(B[55]), .ZN(net446539) );
  NAND2_X1 U357 ( .A1(B[36]), .A2(A[36]), .ZN(n290) );
  NAND2_X1 U358 ( .A1(B[45]), .A2(A[45]), .ZN(n183) );
  NAND2_X1 U360 ( .A1(B[32]), .A2(A[32]), .ZN(n323) );
  OR2_X1 U361 ( .A1(A[27]), .A2(B[27]), .ZN(n380) );
  NAND2_X1 U362 ( .A1(A[42]), .A2(B[42]), .ZN(n216) );
  NAND2_X1 U363 ( .A1(A[40]), .A2(B[40]), .ZN(n265) );
  OR2_X1 U364 ( .A1(B[39]), .A2(A[39]), .ZN(n239) );
  NAND2_X1 U365 ( .A1(A[52]), .A2(B[52]), .ZN(n152) );
  NAND2_X1 U366 ( .A1(B[44]), .A2(A[44]), .ZN(n203) );
  OR2_X1 U367 ( .A1(B[30]), .A2(A[30]), .ZN(n342) );
  NAND2_X1 U368 ( .A1(B[34]), .A2(A[34]), .ZN(n324) );
  OR2_X1 U369 ( .A1(B[26]), .A2(A[26]), .ZN(n385) );
  OR2_X1 U370 ( .A1(B[37]), .A2(A[37]), .ZN(n287) );
  NAND2_X1 U371 ( .A1(B[30]), .A2(A[30]), .ZN(n344) );
  NAND2_X1 U372 ( .A1(B[26]), .A2(A[26]), .ZN(n382) );
  NAND2_X1 U373 ( .A1(B[33]), .A2(A[33]), .ZN(n325) );
  NAND2_X1 U374 ( .A1(B[37]), .A2(A[37]), .ZN(n289) );
  OR2_X1 U375 ( .A1(B[25]), .A2(A[25]), .ZN(n383) );
  NAND2_X1 U376 ( .A1(B[41]), .A2(A[41]), .ZN(n264) );
  NOR2_X1 U377 ( .A1(A[45]), .A2(B[45]), .ZN(n227) );
  NAND2_X1 U378 ( .A1(B[38]), .A2(A[38]), .ZN(n292) );
  NAND2_X1 U379 ( .A1(B[28]), .A2(A[28]), .ZN(n347) );
  OR2_X1 U380 ( .A1(B[28]), .A2(A[28]), .ZN(n359) );
  NAND2_X1 U381 ( .A1(B[29]), .A2(A[29]), .ZN(n345) );
  OR2_X1 U382 ( .A1(B[34]), .A2(A[34]), .ZN(n317) );
  NAND2_X1 U383 ( .A1(B[48]), .A2(A[48]), .ZN(n198) );
  OR2_X1 U384 ( .A1(B[36]), .A2(A[36]), .ZN(n296) );
  OR2_X1 U385 ( .A1(B[21]), .A2(A[21]), .ZN(n408) );
  NAND2_X1 U386 ( .A1(A[27]), .A2(B[27]), .ZN(n381) );
  NAND2_X1 U387 ( .A1(B[31]), .A2(A[31]), .ZN(n338) );
  OR2_X1 U388 ( .A1(A[56]), .A2(B[56]), .ZN(n51) );
  OR2_X1 U389 ( .A1(B[32]), .A2(A[32]), .ZN(n315) );
  OR2_X1 U390 ( .A1(A[29]), .A2(B[29]), .ZN(n360) );
  OR2_X1 U391 ( .A1(B[33]), .A2(A[33]), .ZN(n316) );
  OR2_X1 U392 ( .A1(A[40]), .A2(B[40]), .ZN(n283) );
  OR2_X1 U393 ( .A1(A[31]), .A2(B[31]), .ZN(n343) );
  OR2_X1 U394 ( .A1(A[52]), .A2(B[52]), .ZN(n153) );
  NAND2_X1 U395 ( .A1(B[39]), .A2(A[39]), .ZN(n291) );
  OR2_X1 U396 ( .A1(A[63]), .A2(B[63]), .ZN(n87) );
  OR2_X1 U397 ( .A1(A[62]), .A2(B[62]), .ZN(n93) );
  OR2_X1 U398 ( .A1(A[35]), .A2(B[35]), .ZN(n41) );
  OR2_X1 U399 ( .A1(A[51]), .A2(B[51]), .ZN(n164) );
  AND2_X1 U400 ( .A1(n36), .A2(net446511), .ZN(net537208) );
  AND3_X1 U401 ( .A1(net446505), .A2(n565), .A3(n564), .ZN(n36) );
  INV_X1 U402 ( .A(net446517), .ZN(n564) );
  OR2_X1 U403 ( .A1(B[22]), .A2(A[22]), .ZN(n409) );
  OR2_X1 U404 ( .A1(B[18]), .A2(A[18]), .ZN(n429) );
  OR2_X1 U405 ( .A1(B[14]), .A2(A[14]), .ZN(n462) );
  OR2_X1 U406 ( .A1(B[19]), .A2(A[19]), .ZN(n430) );
  OR2_X1 U407 ( .A1(B[23]), .A2(A[23]), .ZN(n404) );
  OR2_X1 U408 ( .A1(B[16]), .A2(A[16]), .ZN(n437) );
  OR2_X1 U409 ( .A1(B[17]), .A2(A[17]), .ZN(n438) );
  OR2_X1 U410 ( .A1(B[13]), .A2(A[13]), .ZN(n469) );
  OR2_X1 U411 ( .A1(B[20]), .A2(A[20]), .ZN(n412) );
  OR2_X1 U412 ( .A1(B[24]), .A2(A[24]), .ZN(n388) );
  OR2_X1 U413 ( .A1(B[15]), .A2(A[15]), .ZN(n463) );
  OR2_X1 U414 ( .A1(B[6]), .A2(A[6]), .ZN(n78) );
  OR2_X1 U415 ( .A1(B[10]), .A2(A[10]), .ZN(n494) );
  OR2_X1 U416 ( .A1(B[5]), .A2(A[5]), .ZN(n83) );
  OR2_X1 U417 ( .A1(B[9]), .A2(A[9]), .ZN(n65) );
  OR2_X1 U418 ( .A1(B[11]), .A2(A[11]), .ZN(n488) );
  OR2_X1 U419 ( .A1(B[7]), .A2(A[7]), .ZN(n73) );
  OR2_X1 U420 ( .A1(B[8]), .A2(A[8]), .ZN(n69) );
  OR2_X1 U421 ( .A1(B[2]), .A2(A[2]), .ZN(n304) );
  OR2_X1 U422 ( .A1(B[12]), .A2(A[12]), .ZN(n468) );
  OR2_X1 U423 ( .A1(B[1]), .A2(A[1]), .ZN(n372) );
  OR2_X1 U424 ( .A1(B[4]), .A2(A[4]), .ZN(n108) );
  INV_X1 U425 ( .A(B[46]), .ZN(n605) );
  OR2_X1 U426 ( .A1(B[3]), .A2(A[3]), .ZN(n299) );
  OR2_X1 U427 ( .A1(B[0]), .A2(A[0]), .ZN(n508) );
  NAND2_X1 U428 ( .A1(B[1]), .A2(A[1]), .ZN(n371) );
  NAND2_X1 U429 ( .A1(B[8]), .A2(A[8]), .ZN(n70) );
  NAND2_X1 U430 ( .A1(B[12]), .A2(A[12]), .ZN(n459) );
  NAND2_X1 U431 ( .A1(B[14]), .A2(A[14]), .ZN(n461) );
  NAND2_X1 U432 ( .A1(B[24]), .A2(A[24]), .ZN(n387) );
  NAND2_X1 U433 ( .A1(B[17]), .A2(A[17]), .ZN(n434) );
  NAND2_X1 U434 ( .A1(B[4]), .A2(A[4]), .ZN(n107) );
  NAND2_X1 U435 ( .A1(B[13]), .A2(A[13]), .ZN(n460) );
  NAND2_X1 U436 ( .A1(B[22]), .A2(A[22]), .ZN(n406) );
  NAND2_X1 U437 ( .A1(B[16]), .A2(A[16]), .ZN(n436) );
  NAND2_X1 U438 ( .A1(B[25]), .A2(A[25]), .ZN(n386) );
  NAND2_X1 U439 ( .A1(B[5]), .A2(A[5]), .ZN(n82) );
  NAND2_X1 U440 ( .A1(B[9]), .A2(A[9]), .ZN(n66) );
  NAND2_X1 U441 ( .A1(B[18]), .A2(A[18]), .ZN(n433) );
  NAND2_X1 U442 ( .A1(B[2]), .A2(A[2]), .ZN(n301) );
  NAND2_X1 U443 ( .A1(B[0]), .A2(A[0]), .ZN(n441) );
  NAND2_X1 U444 ( .A1(B[6]), .A2(A[6]), .ZN(n75) );
  NAND2_X1 U445 ( .A1(B[10]), .A2(A[10]), .ZN(n491) );
  NAND2_X1 U446 ( .A1(B[21]), .A2(A[21]), .ZN(n410) );
  NAND2_X1 U447 ( .A1(B[20]), .A2(A[20]), .ZN(n411) );
  NAND2_X1 U448 ( .A1(B[3]), .A2(A[3]), .ZN(n300) );
  NAND2_X1 U449 ( .A1(B[15]), .A2(A[15]), .ZN(n457) );
  NAND2_X1 U450 ( .A1(B[19]), .A2(A[19]), .ZN(n428) );
  NAND2_X1 U451 ( .A1(B[23]), .A2(A[23]), .ZN(n405) );
  NAND2_X1 U452 ( .A1(B[7]), .A2(A[7]), .ZN(n74) );
  NAND2_X1 U453 ( .A1(B[11]), .A2(A[11]), .ZN(n492) );
  XNOR2_X1 U454 ( .A(n242), .B(n241), .ZN(SUM[47]) );
  OR2_X1 U455 ( .A1(A[59]), .A2(B[59]), .ZN(net446522) );
  NAND4_X1 U456 ( .A1(n161), .A2(n162), .A3(n193), .A4(n163), .ZN(n160) );
  INV_X1 U457 ( .A(n163), .ZN(n576) );
  OAI211_X1 U458 ( .C1(n575), .C2(n174), .A(n163), .B(n175), .ZN(n172) );
  OAI21_X1 U459 ( .B1(n61), .B2(n101), .A(net446539), .ZN(n119) );
  NOR2_X1 U460 ( .A1(n572), .A2(n125), .ZN(n117) );
  NAND2_X1 U461 ( .A1(A[47]), .A2(B[47]), .ZN(n180) );
  OR2_X1 U462 ( .A1(A[47]), .A2(B[47]), .ZN(n211) );
  OR2_X1 U463 ( .A1(A[47]), .A2(B[47]), .ZN(n6) );
  XNOR2_X1 U464 ( .A(n25), .B(n252), .ZN(SUM[45]) );
  NAND2_X1 U465 ( .A1(A[43]), .A2(B[43]), .ZN(n215) );
  AOI211_X1 U466 ( .C1(n127), .C2(n128), .A(net446593), .B(n129), .ZN(n126) );
  NAND4_X1 U467 ( .A1(n231), .A2(n228), .A3(n230), .A4(n28), .ZN(n177) );
  INV_X1 U468 ( .A(n230), .ZN(n552) );
  NOR2_X1 U469 ( .A1(n132), .A2(n125), .ZN(n128) );
  INV_X1 U470 ( .A(net446521), .ZN(n563) );
  NAND2_X1 U471 ( .A1(n51), .A2(net446521), .ZN(n115) );
  AOI21_X1 U472 ( .B1(n566), .B2(net446521), .A(n562), .ZN(n116) );
  NAND2_X1 U473 ( .A1(A[49]), .A2(B[49]), .ZN(n193) );
  OR2_X2 U474 ( .A1(A[57]), .A2(B[57]), .ZN(net446521) );
  AOI21_X1 U475 ( .B1(n14), .B2(n27), .A(n148), .ZN(n149) );
  AND2_X1 U476 ( .A1(n164), .A2(n123), .ZN(n4) );
  NAND4_X1 U477 ( .A1(n164), .A2(n166), .A3(n165), .A4(n167), .ZN(n122) );
  AND2_X1 U478 ( .A1(n164), .A2(n165), .ZN(n159) );
  XNOR2_X1 U479 ( .A(n534), .B(n309), .ZN(SUM[38]) );
  NAND2_X1 U480 ( .A1(n534), .A2(n237), .ZN(n307) );
  NOR2_X1 U481 ( .A1(net446512), .A2(net537208), .ZN(net446509) );
  OAI21_X1 U482 ( .B1(n130), .B2(n61), .A(net446534), .ZN(n129) );
  INV_X1 U483 ( .A(net446516), .ZN(n570) );
  OAI21_X1 U484 ( .B1(n217), .B2(n541), .A(n219), .ZN(n213) );
  NAND2_X1 U485 ( .A1(n50), .A2(n103), .ZN(n112) );
  NAND2_X1 U486 ( .A1(net446519), .A2(n50), .ZN(n130) );
  NAND2_X1 U487 ( .A1(A[59]), .A2(B[59]), .ZN(net446516) );
  XNOR2_X1 U488 ( .A(n169), .B(n4), .ZN(SUM[51]) );
  AOI21_X1 U489 ( .B1(n280), .B2(n281), .A(n548), .ZN(n279) );
  NAND2_X1 U490 ( .A1(n285), .A2(n286), .ZN(n281) );
  XNOR2_X1 U491 ( .A(n272), .B(n274), .ZN(SUM[42]) );
  NAND2_X1 U492 ( .A1(n10), .A2(n133), .ZN(n101) );
  INV_X1 U493 ( .A(n133), .ZN(n572) );
  NAND2_X1 U494 ( .A1(B[53]), .A2(A[53]), .ZN(n121) );
  AND2_X1 U495 ( .A1(n141), .A2(n140), .ZN(n50) );
  OR2_X1 U496 ( .A1(A[54]), .A2(B[54]), .ZN(n140) );
  OR2_X1 U497 ( .A1(A[55]), .A2(B[55]), .ZN(n141) );
  NAND2_X1 U498 ( .A1(n605), .A2(n553), .ZN(n230) );
  NAND2_X1 U499 ( .A1(B[58]), .A2(A[58]), .ZN(net446535) );
  XNOR2_X1 U500 ( .A(n329), .B(n330), .ZN(SUM[34]) );
  NAND2_X1 U501 ( .A1(n317), .A2(n329), .ZN(n328) );
  NAND4_X1 U502 ( .A1(n335), .A2(n336), .A3(n337), .A4(n338), .ZN(n28) );
  NAND4_X1 U503 ( .A1(n335), .A2(n336), .A3(n337), .A4(n338), .ZN(n229) );
  XNOR2_X1 U504 ( .A(n94), .B(n95), .ZN(SUM[63]) );
  AOI21_X1 U505 ( .B1(n117), .B2(n118), .A(n119), .ZN(n114) );
  AOI21_X1 U506 ( .B1(n118), .B2(n153), .A(n559), .ZN(n154) );
  OAI211_X1 U507 ( .C1(net538658), .C2(n569), .A(net446490), .B(net446491), 
        .ZN(net446484) );
  NAND2_X1 U508 ( .A1(n90), .A2(n87), .ZN(n94) );
  OAI211_X1 U509 ( .C1(n563), .C2(net446534), .A(net446535), .B(n515), .ZN(n38) );
  AND2_X1 U510 ( .A1(net446536), .A2(net446521), .ZN(net446587) );
  AND3_X1 U511 ( .A1(net446536), .A2(net446539), .A3(net446534), .ZN(net535419) );
  INV_X1 U512 ( .A(net446536), .ZN(n562) );
  NAND2_X1 U513 ( .A1(n321), .A2(n519), .ZN(n327) );
  NAND4_X1 U514 ( .A1(n41), .A2(n54), .A3(n317), .A4(n28), .ZN(n314) );
  NAND2_X1 U515 ( .A1(n159), .A2(n160), .ZN(n124) );
  XNOR2_X1 U516 ( .A(n269), .B(n270), .ZN(SUM[43]) );
  NAND2_X1 U517 ( .A1(B[63]), .A2(A[63]), .ZN(n90) );
  NOR2_X1 U518 ( .A1(n62), .A2(n145), .ZN(n144) );
  NOR2_X1 U519 ( .A1(B[53]), .A2(A[53]), .ZN(n138) );
  XNOR2_X1 U520 ( .A(net446508), .B(net446509), .ZN(SUM[61]) );
  NAND2_X1 U521 ( .A1(A[57]), .A2(B[57]), .ZN(net446536) );
  NAND2_X1 U524 ( .A1(n257), .A2(n520), .ZN(n260) );
  AND3_X1 U525 ( .A1(n6), .A2(n234), .A3(n520), .ZN(n208) );
  AND2_X1 U526 ( .A1(n263), .A2(n256), .ZN(n9) );
  INV_X1 U527 ( .A(n256), .ZN(n545) );
  AND2_X1 U530 ( .A1(n263), .A2(n256), .ZN(n268) );
  NAND2_X1 U533 ( .A1(net446520), .A2(net446521), .ZN(n104) );
  AND2_X1 U534 ( .A1(net446522), .A2(net446520), .ZN(n37) );
  NAND2_X1 U535 ( .A1(net446520), .A2(net446535), .ZN(net446564) );
  OAI211_X1 U536 ( .C1(A[59]), .C2(B[59]), .A(net446520), .B(net446521), .ZN(
        net446517) );
  OAI211_X1 U537 ( .C1(n562), .C2(n51), .A(net446521), .B(net446520), .ZN(n35)
         );
  OAI211_X1 U538 ( .C1(n122), .C2(n52), .A(n518), .B(n123), .ZN(n118) );
  OAI211_X1 U539 ( .C1(n52), .C2(n122), .A(n123), .B(n124), .ZN(n127) );
  OAI211_X1 U540 ( .C1(n52), .C2(n122), .A(n123), .B(n518), .ZN(n27) );
  XNOR2_X1 U541 ( .A(n144), .B(n57), .ZN(SUM[55]) );
  OR2_X1 U542 ( .A1(B[50]), .A2(A[50]), .ZN(n165) );
  NAND2_X1 U545 ( .A1(A[50]), .A2(B[50]), .ZN(n163) );
  NAND2_X1 U546 ( .A1(net446513), .A2(net446516), .ZN(net446530) );
  NAND2_X1 U547 ( .A1(n37), .A2(n38), .ZN(net446513) );
  XNOR2_X1 U548 ( .A(n92), .B(net446526), .ZN(SUM[60]) );
  AOI21_X1 U549 ( .B1(n99), .B2(net446511), .A(net446530), .ZN(n92) );
  AND2_X1 U550 ( .A1(n93), .A2(net538437), .ZN(n88) );
  NAND2_X1 U552 ( .A1(net538437), .A2(net446505), .ZN(net446501) );
  AND2_X1 U554 ( .A1(net538437), .A2(net446490), .ZN(net446508) );
  INV_X1 U555 ( .A(n30), .ZN(n534) );
  OAI21_X1 U556 ( .B1(B[35]), .B2(A[35]), .A(n317), .ZN(n31) );
  NAND2_X1 U557 ( .A1(A[35]), .A2(B[35]), .ZN(n321) );
  NAND2_X1 U559 ( .A1(B[54]), .A2(A[54]), .ZN(n131) );
  XNOR2_X1 U563 ( .A(n113), .B(net446564), .ZN(SUM[58]) );
  NAND2_X1 U564 ( .A1(n90), .A2(n91), .ZN(n89) );
  NAND2_X1 U565 ( .A1(n91), .A2(n96), .ZN(n95) );
  NAND2_X1 U566 ( .A1(n93), .A2(n91), .ZN(n98) );
  XNOR2_X1 U567 ( .A(n158), .B(n127), .ZN(SUM[52]) );
  XNOR2_X1 U568 ( .A(n126), .B(net446587), .ZN(SUM[57]) );
  NOR2_X1 U569 ( .A1(B[56]), .A2(A[56]), .ZN(net446594) );
  NAND2_X1 U570 ( .A1(A[56]), .A2(B[56]), .ZN(net446534) );
  OR2_X1 U571 ( .A1(A[56]), .A2(B[56]), .ZN(net446519) );
  NOR2_X1 U572 ( .A1(A[46]), .A2(B[46]), .ZN(n226) );
  NAND2_X1 U573 ( .A1(B[46]), .A2(A[46]), .ZN(n185) );
  INV_X1 U576 ( .A(A[46]), .ZN(n553) );
  OAI21_X1 U577 ( .B1(n114), .B2(n115), .A(n116), .ZN(n113) );
  NAND2_X1 U578 ( .A1(B[62]), .A2(A[62]), .ZN(n91) );
  NOR2_X1 U579 ( .A1(n138), .A2(n137), .ZN(n135) );
  OAI21_X1 U580 ( .B1(n152), .B2(n138), .A(n121), .ZN(n148) );
  AOI21_X1 U581 ( .B1(n561), .B2(n111), .A(n571), .ZN(n109) );
  INV_X1 U582 ( .A(n35), .ZN(n561) );
  AND2_X1 U583 ( .A1(net446522), .A2(net446516), .ZN(net537284) );
  XNOR2_X1 U584 ( .A(n149), .B(n150), .ZN(SUM[54]) );
  NAND2_X1 U585 ( .A1(A[51]), .A2(B[51]), .ZN(n123) );
  NAND2_X1 U586 ( .A1(n224), .A2(n314), .ZN(n45) );
  OAI211_X1 U587 ( .C1(n31), .C2(n537), .A(n321), .B(n314), .ZN(n293) );
  NAND2_X1 U588 ( .A1(B[61]), .A2(A[61]), .ZN(net446490) );
  NAND4_X1 U589 ( .A1(n27), .A2(n135), .A3(n10), .A4(n133), .ZN(n102) );
  NAND2_X1 U590 ( .A1(n133), .A2(n51), .ZN(n132) );
  NAND2_X1 U591 ( .A1(n148), .A2(n140), .ZN(n146) );
  INV_X1 U592 ( .A(net446490), .ZN(n568) );
  OAI21_X1 U593 ( .B1(net538658), .B2(net446501), .A(net446502), .ZN(n97) );
  AOI21_X1 U594 ( .B1(n526), .B2(net538437), .A(n568), .ZN(net446502) );
  NOR2_X1 U595 ( .A1(n526), .A2(n569), .ZN(net446526) );
  OAI21_X1 U596 ( .B1(net446513), .B2(n569), .A(net446514), .ZN(net446512) );
  XNOR2_X1 U597 ( .A(n97), .B(n98), .ZN(SUM[62]) );
  NAND2_X1 U598 ( .A1(n93), .A2(n97), .ZN(n96) );
  AOI21_X1 U599 ( .B1(n570), .B2(net446505), .A(n526), .ZN(net446514) );
endmodule


module RCA_NBIT64_3 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_3_DW01_add_5 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_2_DW01_add_3 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net431092, net431087, net431086, net431073, net431072, net431070,
         net431069, net431061, net431059, net431057, net537977, net538409,
         net431081, net431068, net431076, net431065, net431064, n1, n2, n3, n4,
         n5, n8, n10, n11, n12, n14, n15, n16, n20, n21, n23, n24, n28, n29,
         n30, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n46, n47, n51,
         n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n68, n69,
         n70, n71, n72, n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n109, n110, n111, n112, n113,
         n114, n115, n116, n118, n119, n120, n121, n123, n125, n126, n127,
         n129, n130, n131, n132, n133, n134, n135, n136, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n164, n165,
         n166, n167, n168, n169, n170, n172, n174, n176, n177, n178, n179,
         n180, n181, n182, n183, n185, n186, n187, n188, n189, n190, n191,
         n193, n194, n195, n196, n197, n198, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n215, n216, n218,
         n219, n220, n222, n224, n226, n227, n230, n231, n232, n233, n234,
         n235, n236, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n260, n261, n262, n263, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n292, n293, n294, n295,
         n296, n297, n298, n299, n301, n302, n303, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n332, n334, n335, n336, n339, n340, n341, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n354, n356, n357, n358, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n377, n378, n380, n381, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n402, n404, n405, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n429, n430, n431, n432, n433, n434, n435,
         n436, n438, n440, n441, n442, n443, n444, n447, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n483, n484, n485, n486, n489,
         n490, n491, n492, n493, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575;

  NAND3_X1 U42 ( .A1(n28), .A2(n183), .A3(n182), .ZN(n29) );
  OR2_X2 U53 ( .A1(B[52]), .A2(A[52]), .ZN(n153) );
  NAND3_X1 U59 ( .A1(n46), .A2(n183), .A3(n182), .ZN(n150) );
  NAND3_X1 U60 ( .A1(net431070), .A2(net431069), .A3(net431065), .ZN(n35) );
  NAND3_X1 U520 ( .A1(n29), .A2(n149), .A3(n148), .ZN(n147) );
  NAND3_X1 U534 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n244) );
  NAND3_X1 U535 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n245) );
  NAND3_X1 U575 ( .A1(n471), .A2(n472), .A3(n473), .ZN(n470) );
  NAND3_X1 U576 ( .A1(n474), .A2(n78), .A3(n475), .ZN(n471) );
  NAND3_X1 U581 ( .A1(n485), .A2(n88), .A3(n87), .ZN(n484) );
  NAND3_X1 U582 ( .A1(n96), .A2(n486), .A3(n91), .ZN(n485) );
  CLKBUF_X1 U2 ( .A(n47), .Z(n496) );
  AND2_X1 U3 ( .A1(n489), .A2(n422), .ZN(SUM[0]) );
  OR2_X1 U4 ( .A1(A[60]), .A2(B[60]), .ZN(net431069) );
  CLKBUF_X1 U5 ( .A(A[47]), .Z(n497) );
  OR2_X1 U6 ( .A1(B[57]), .A2(A[57]), .ZN(n114) );
  CLKBUF_X1 U7 ( .A(A[59]), .Z(n498) );
  CLKBUF_X1 U8 ( .A(n253), .Z(n499) );
  CLKBUF_X1 U9 ( .A(n57), .Z(n500) );
  AND2_X1 U10 ( .A1(n21), .A2(n11), .ZN(n501) );
  XNOR2_X1 U11 ( .A(n164), .B(n502), .ZN(SUM[55]) );
  AND2_X1 U12 ( .A1(n539), .A2(n156), .ZN(n502) );
  CLKBUF_X1 U13 ( .A(n24), .Z(n504) );
  CLKBUF_X1 U14 ( .A(A[51]), .Z(n503) );
  NOR2_X1 U15 ( .A1(A[49]), .A2(B[49]), .ZN(n54) );
  OR2_X1 U16 ( .A1(B[53]), .A2(A[53]), .ZN(n155) );
  OR2_X2 U17 ( .A1(A[42]), .A2(B[42]), .ZN(n250) );
  AND4_X2 U18 ( .A1(n254), .A2(n248), .A3(n250), .A4(n243), .ZN(n21) );
  NOR2_X1 U19 ( .A1(A[51]), .A2(B[51]), .ZN(n505) );
  NOR2_X1 U20 ( .A1(B[50]), .A2(A[50]), .ZN(n57) );
  AND3_X1 U21 ( .A1(n226), .A2(n213), .A3(n507), .ZN(n506) );
  AND2_X1 U22 ( .A1(n215), .A2(n227), .ZN(n507) );
  AND3_X1 U23 ( .A1(n226), .A2(n213), .A3(n507), .ZN(n59) );
  NAND2_X1 U24 ( .A1(n506), .A2(n501), .ZN(n205) );
  OR2_X2 U25 ( .A1(A[45]), .A2(B[45]), .ZN(n215) );
  XOR2_X1 U26 ( .A(n239), .B(n508), .Z(SUM[45]) );
  NAND2_X1 U27 ( .A1(n63), .A2(n64), .ZN(n508) );
  INV_X1 U28 ( .A(n380), .ZN(n551) );
  INV_X1 U29 ( .A(n420), .ZN(n560) );
  INV_X1 U30 ( .A(n35), .ZN(n515) );
  OAI21_X1 U31 ( .B1(n573), .B2(n456), .A(n453), .ZN(n81) );
  OAI21_X1 U32 ( .B1(n560), .B2(n341), .A(n556), .ZN(n394) );
  INV_X1 U33 ( .A(n332), .ZN(n556) );
  OAI21_X1 U34 ( .B1(n555), .B2(n335), .A(n334), .ZN(n380) );
  INV_X1 U35 ( .A(n394), .ZN(n555) );
  OAI21_X1 U36 ( .B1(n551), .B2(n329), .A(n330), .ZN(n357) );
  AOI21_X1 U37 ( .B1(n452), .B2(n453), .A(n454), .ZN(n447) );
  NAND2_X1 U38 ( .A1(n568), .A2(n455), .ZN(n452) );
  INV_X1 U39 ( .A(n456), .ZN(n568) );
  OAI21_X1 U40 ( .B1(n328), .B2(n329), .A(n330), .ZN(n327) );
  AOI21_X1 U41 ( .B1(n550), .B2(n332), .A(n552), .ZN(n328) );
  INV_X1 U43 ( .A(n334), .ZN(n552) );
  INV_X1 U44 ( .A(n335), .ZN(n550) );
  NAND2_X1 U45 ( .A1(n433), .A2(n434), .ZN(n420) );
  OAI21_X1 U46 ( .B1(n447), .B2(n565), .A(n14), .ZN(n433) );
  AOI21_X1 U47 ( .B1(n435), .B2(n436), .A(n561), .ZN(n434) );
  INV_X1 U48 ( .A(n451), .ZN(n565) );
  NOR2_X1 U49 ( .A1(n560), .A2(n335), .ZN(n336) );
  NAND2_X1 U50 ( .A1(n468), .A2(n451), .ZN(n466) );
  NAND2_X1 U51 ( .A1(n564), .A2(n81), .ZN(n468) );
  INV_X1 U52 ( .A(n454), .ZN(n564) );
  INV_X1 U54 ( .A(n455), .ZN(n573) );
  INV_X1 U55 ( .A(n329), .ZN(n546) );
  INV_X1 U56 ( .A(n341), .ZN(n557) );
  INV_X1 U57 ( .A(n98), .ZN(SUM[64]) );
  NOR2_X1 U58 ( .A1(n540), .A2(n541), .ZN(n136) );
  INV_X1 U61 ( .A(n119), .ZN(n540) );
  AND2_X1 U62 ( .A1(n120), .A2(n71), .ZN(n1) );
  NAND2_X1 U63 ( .A1(n208), .A2(n210), .ZN(n232) );
  NAND2_X1 U64 ( .A1(n269), .A2(n288), .ZN(n287) );
  NAND2_X1 U65 ( .A1(n139), .A2(n113), .ZN(n144) );
  NAND2_X1 U66 ( .A1(n191), .A2(n543), .ZN(n196) );
  INV_X1 U67 ( .A(n139), .ZN(n532) );
  XNOR2_X1 U68 ( .A(n169), .B(n170), .ZN(SUM[54]) );
  NOR2_X1 U69 ( .A1(n536), .A2(n73), .ZN(n170) );
  AOI21_X1 U70 ( .B1(n172), .B2(n155), .A(n542), .ZN(n169) );
  INV_X1 U71 ( .A(n161), .ZN(n536) );
  NAND2_X1 U72 ( .A1(n155), .A2(n159), .ZN(n177) );
  NAND2_X1 U73 ( .A1(n273), .A2(n269), .ZN(n290) );
  NAND2_X1 U74 ( .A1(n168), .A2(n153), .ZN(n180) );
  NAND2_X1 U75 ( .A1(n254), .A2(n252), .ZN(n263) );
  NAND4_X1 U76 ( .A1(n317), .A2(n318), .A3(n319), .A4(n320), .ZN(n230) );
  NAND2_X1 U77 ( .A1(n72), .A2(n327), .ZN(n318) );
  NAND4_X1 U78 ( .A1(n336), .A2(n557), .A3(n546), .A4(n72), .ZN(n317) );
  NAND2_X1 U79 ( .A1(n2), .A2(n326), .ZN(n319) );
  OAI21_X1 U80 ( .B1(n4), .B2(n518), .A(n306), .ZN(n311) );
  AND2_X1 U81 ( .A1(n315), .A2(n305), .ZN(n4) );
  OAI21_X1 U82 ( .B1(n348), .B2(n3), .A(n323), .ZN(n346) );
  XNOR2_X1 U83 ( .A(n230), .B(n316), .ZN(SUM[32]) );
  NAND2_X1 U84 ( .A1(n296), .A2(n305), .ZN(n316) );
  OAI21_X1 U85 ( .B1(n516), .B2(n231), .A(n224), .ZN(n253) );
  INV_X1 U86 ( .A(n277), .ZN(n516) );
  XNOR2_X1 U87 ( .A(net538409), .B(net431092), .ZN(SUM[60]) );
  NAND2_X1 U88 ( .A1(net431068), .A2(net431069), .ZN(net431092) );
  XNOR2_X1 U89 ( .A(n295), .B(n277), .ZN(SUM[36]) );
  NAND2_X1 U90 ( .A1(n276), .A2(n275), .ZN(n295) );
  XNOR2_X1 U91 ( .A(n311), .B(n312), .ZN(SUM[34]) );
  NAND2_X1 U92 ( .A1(n298), .A2(n307), .ZN(n312) );
  XNOR2_X1 U93 ( .A(n43), .B(n236), .ZN(SUM[46]) );
  NAND2_X1 U94 ( .A1(n213), .A2(n524), .ZN(n236) );
  OAI21_X1 U95 ( .B1(n58), .B2(n523), .A(n212), .ZN(n43) );
  XNOR2_X1 U96 ( .A(n313), .B(n314), .ZN(SUM[33]) );
  NAND2_X1 U97 ( .A1(n315), .A2(n305), .ZN(n313) );
  NAND2_X1 U98 ( .A1(n297), .A2(n306), .ZN(n314) );
  XNOR2_X1 U99 ( .A(n343), .B(n344), .ZN(SUM[31]) );
  NAND2_X1 U100 ( .A1(n320), .A2(n326), .ZN(n343) );
  NAND2_X1 U101 ( .A1(n324), .A2(n345), .ZN(n344) );
  NAND2_X1 U102 ( .A1(n346), .A2(n325), .ZN(n345) );
  XNOR2_X1 U103 ( .A(n202), .B(n203), .ZN(SUM[49]) );
  NAND2_X1 U104 ( .A1(n190), .A2(n544), .ZN(n202) );
  XNOR2_X1 U105 ( .A(n241), .B(n240), .ZN(SUM[44]) );
  NAND2_X1 U106 ( .A1(n227), .A2(n216), .ZN(n241) );
  XNOR2_X1 U107 ( .A(n260), .B(n261), .ZN(SUM[41]) );
  NAND2_X1 U108 ( .A1(n248), .A2(n251), .ZN(n261) );
  NAND2_X1 U109 ( .A1(n262), .A2(n252), .ZN(n260) );
  XNOR2_X1 U110 ( .A(n5), .B(n258), .ZN(SUM[42]) );
  NAND2_X1 U111 ( .A1(n250), .A2(n246), .ZN(n258) );
  OAI21_X1 U112 ( .B1(n51), .B2(n527), .A(n251), .ZN(n5) );
  XNOR2_X1 U113 ( .A(n293), .B(n292), .ZN(SUM[37]) );
  NAND2_X1 U114 ( .A1(n271), .A2(n274), .ZN(n293) );
  NAND2_X1 U115 ( .A1(n294), .A2(n275), .ZN(n292) );
  XNOR2_X1 U116 ( .A(n346), .B(n347), .ZN(SUM[30]) );
  NAND2_X1 U117 ( .A1(n325), .A2(n324), .ZN(n347) );
  XNOR2_X1 U118 ( .A(n370), .B(n371), .ZN(SUM[27]) );
  NAND2_X1 U119 ( .A1(n363), .A2(n372), .ZN(n370) );
  NAND2_X1 U120 ( .A1(n361), .A2(n362), .ZN(n371) );
  NAND2_X1 U121 ( .A1(n373), .A2(n366), .ZN(n372) );
  XNOR2_X1 U122 ( .A(n348), .B(n354), .ZN(SUM[29]) );
  NOR2_X1 U123 ( .A1(n545), .A2(n3), .ZN(n354) );
  INV_X1 U124 ( .A(n323), .ZN(n545) );
  NAND2_X1 U125 ( .A1(n215), .A2(n212), .ZN(n239) );
  XNOR2_X1 U126 ( .A(n358), .B(n357), .ZN(SUM[28]) );
  NAND2_X1 U127 ( .A1(n339), .A2(n322), .ZN(n358) );
  XNOR2_X1 U128 ( .A(n378), .B(n377), .ZN(SUM[25]) );
  NAND2_X1 U129 ( .A1(n364), .A2(n367), .ZN(n378) );
  XNOR2_X1 U130 ( .A(n374), .B(n373), .ZN(SUM[26]) );
  NAND2_X1 U131 ( .A1(n366), .A2(n363), .ZN(n374) );
  OAI21_X1 U132 ( .B1(n517), .B2(n301), .A(n302), .ZN(n222) );
  INV_X1 U133 ( .A(n303), .ZN(n517) );
  NAND2_X1 U134 ( .A1(n299), .A2(n298), .ZN(n301) );
  OAI211_X1 U135 ( .C1(n518), .C2(n305), .A(n306), .B(n307), .ZN(n303) );
  OAI211_X1 U136 ( .C1(n197), .C2(n54), .A(n190), .B(n198), .ZN(n24) );
  NAND2_X1 U137 ( .A1(n528), .A2(n544), .ZN(n198) );
  XNOR2_X1 U138 ( .A(n308), .B(n309), .ZN(SUM[35]) );
  NAND2_X1 U139 ( .A1(n302), .A2(n299), .ZN(n309) );
  NAND2_X1 U140 ( .A1(n310), .A2(n307), .ZN(n308) );
  NAND2_X1 U141 ( .A1(n311), .A2(n298), .ZN(n310) );
  AOI21_X1 U142 ( .B1(n10), .B2(n512), .A(n73), .ZN(n164) );
  AND2_X1 U143 ( .A1(n155), .A2(n161), .ZN(n10) );
  OAI21_X1 U144 ( .B1(n20), .B2(n519), .A(n274), .ZN(n289) );
  INV_X1 U145 ( .A(n271), .ZN(n519) );
  AND2_X1 U146 ( .A1(n294), .A2(n275), .ZN(n20) );
  AND2_X1 U147 ( .A1(n148), .A2(n149), .ZN(n181) );
  NAND4_X1 U148 ( .A1(n267), .A2(n271), .A3(n273), .A4(n276), .ZN(n231) );
  XNOR2_X1 U149 ( .A(n256), .B(n255), .ZN(SUM[43]) );
  NAND2_X1 U150 ( .A1(n257), .A2(n246), .ZN(n256) );
  NAND2_X1 U151 ( .A1(n251), .A2(n252), .ZN(n249) );
  OR2_X1 U152 ( .A1(n69), .A2(n222), .ZN(n277) );
  AND2_X1 U153 ( .A1(n70), .A2(n230), .ZN(n69) );
  AND4_X1 U154 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n70) );
  NOR2_X1 U155 ( .A1(n54), .A2(n529), .ZN(n182) );
  INV_X1 U156 ( .A(n185), .ZN(n529) );
  NOR2_X1 U157 ( .A1(n509), .A2(n510), .ZN(n11) );
  NAND2_X1 U158 ( .A1(n522), .A2(n230), .ZN(n509) );
  NAND4_X1 U159 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n510) );
  XNOR2_X1 U160 ( .A(n400), .B(n402), .ZN(SUM[21]) );
  NOR2_X1 U161 ( .A1(n554), .A2(n553), .ZN(n402) );
  INV_X1 U162 ( .A(n391), .ZN(n554) );
  OAI21_X1 U163 ( .B1(n58), .B2(n523), .A(n212), .ZN(n235) );
  OAI21_X1 U164 ( .B1(n51), .B2(n527), .A(n251), .ZN(n23) );
  NAND2_X1 U165 ( .A1(n230), .A2(n296), .ZN(n315) );
  OAI211_X1 U166 ( .C1(n106), .C2(n538), .A(n42), .B(n539), .ZN(n105) );
  NAND2_X1 U167 ( .A1(n161), .A2(n66), .ZN(n106) );
  AND2_X1 U168 ( .A1(n356), .A2(n322), .ZN(n348) );
  NAND2_X1 U169 ( .A1(n357), .A2(n339), .ZN(n356) );
  AND2_X1 U170 ( .A1(n262), .A2(n252), .ZN(n51) );
  NAND2_X1 U171 ( .A1(n277), .A2(n276), .ZN(n294) );
  INV_X1 U172 ( .A(n54), .ZN(n544) );
  INV_X1 U173 ( .A(n215), .ZN(n523) );
  INV_X1 U174 ( .A(n248), .ZN(n527) );
  INV_X1 U175 ( .A(n389), .ZN(n553) );
  NAND2_X1 U176 ( .A1(n159), .A2(n168), .ZN(n167) );
  INV_X1 U177 ( .A(n297), .ZN(n518) );
  NAND2_X1 U178 ( .A1(n174), .A2(n168), .ZN(n172) );
  OAI21_X1 U179 ( .B1(n511), .B2(n176), .A(n153), .ZN(n174) );
  NAND2_X1 U180 ( .A1(n148), .A2(n149), .ZN(n176) );
  INV_X1 U181 ( .A(n159), .ZN(n542) );
  NAND2_X1 U182 ( .A1(n59), .A2(n218), .ZN(n206) );
  AOI21_X1 U183 ( .B1(n522), .B2(n222), .A(n520), .ZN(n219) );
  INV_X1 U184 ( .A(n21), .ZN(n525) );
  NAND2_X1 U185 ( .A1(n153), .A2(n154), .ZN(n152) );
  NAND2_X1 U186 ( .A1(n274), .A2(n275), .ZN(n272) );
  INV_X1 U187 ( .A(n112), .ZN(n541) );
  INV_X1 U188 ( .A(n500), .ZN(n543) );
  INV_X1 U189 ( .A(n216), .ZN(n526) );
  INV_X1 U190 ( .A(n30), .ZN(n539) );
  INV_X1 U191 ( .A(n33), .ZN(n524) );
  AND2_X1 U192 ( .A1(n161), .A2(n66), .ZN(n60) );
  AND2_X1 U193 ( .A1(n121), .A2(n119), .ZN(n71) );
  NAND2_X1 U194 ( .A1(n133), .A2(n119), .ZN(n132) );
  OR2_X1 U195 ( .A1(n526), .A2(n227), .ZN(n64) );
  AND2_X1 U196 ( .A1(n321), .A2(n325), .ZN(n2) );
  OAI211_X1 U197 ( .C1(n3), .C2(n322), .A(n323), .B(n324), .ZN(n321) );
  AND2_X1 U198 ( .A1(n113), .A2(n114), .ZN(n61) );
  XNOR2_X1 U199 ( .A(n423), .B(n424), .ZN(SUM[19]) );
  NAND2_X1 U200 ( .A1(n414), .A2(n425), .ZN(n423) );
  NAND2_X1 U201 ( .A1(n409), .A2(n411), .ZN(n424) );
  NAND2_X1 U202 ( .A1(n426), .A2(n410), .ZN(n425) );
  XNOR2_X1 U203 ( .A(n457), .B(n458), .ZN(SUM[15]) );
  NAND2_X1 U204 ( .A1(n459), .A2(n442), .ZN(n458) );
  NAND2_X1 U205 ( .A1(n438), .A2(n444), .ZN(n457) );
  NAND2_X1 U206 ( .A1(n443), .A2(n460), .ZN(n459) );
  XNOR2_X1 U207 ( .A(n395), .B(n396), .ZN(SUM[23]) );
  NAND2_X1 U208 ( .A1(n387), .A2(n397), .ZN(n396) );
  NAND2_X1 U209 ( .A1(n386), .A2(n385), .ZN(n395) );
  NAND2_X1 U210 ( .A1(n390), .A2(n398), .ZN(n397) );
  XNOR2_X1 U211 ( .A(n432), .B(n420), .ZN(SUM[16]) );
  NAND2_X1 U212 ( .A1(n417), .A2(n418), .ZN(n432) );
  XNOR2_X1 U213 ( .A(n430), .B(n429), .ZN(SUM[17]) );
  NAND2_X1 U214 ( .A1(n419), .A2(n415), .ZN(n430) );
  XNOR2_X1 U215 ( .A(n405), .B(n394), .ZN(SUM[20]) );
  NAND2_X1 U216 ( .A1(n393), .A2(n392), .ZN(n405) );
  XNOR2_X1 U217 ( .A(n381), .B(n380), .ZN(SUM[24]) );
  NAND2_X1 U218 ( .A1(n369), .A2(n368), .ZN(n381) );
  XNOR2_X1 U219 ( .A(n461), .B(n460), .ZN(SUM[14]) );
  NAND2_X1 U220 ( .A1(n443), .A2(n442), .ZN(n461) );
  XNOR2_X1 U221 ( .A(n427), .B(n426), .ZN(SUM[18]) );
  NAND2_X1 U222 ( .A1(n410), .A2(n414), .ZN(n427) );
  XNOR2_X1 U223 ( .A(n399), .B(n398), .ZN(SUM[22]) );
  NAND2_X1 U224 ( .A1(n390), .A2(n387), .ZN(n399) );
  XNOR2_X1 U225 ( .A(n464), .B(n463), .ZN(SUM[13]) );
  NAND2_X1 U226 ( .A1(n450), .A2(n441), .ZN(n464) );
  XNOR2_X1 U227 ( .A(n84), .B(n85), .ZN(SUM[7]) );
  NAND2_X1 U228 ( .A1(n88), .A2(n89), .ZN(n84) );
  NAND2_X1 U229 ( .A1(n86), .A2(n87), .ZN(n85) );
  NAND2_X1 U230 ( .A1(n90), .A2(n91), .ZN(n89) );
  XNOR2_X1 U231 ( .A(n278), .B(n279), .ZN(SUM[3]) );
  NAND2_X1 U232 ( .A1(n282), .A2(n283), .ZN(n278) );
  NAND2_X1 U233 ( .A1(n280), .A2(n281), .ZN(n279) );
  NAND2_X1 U234 ( .A1(n284), .A2(n285), .ZN(n283) );
  XNOR2_X1 U235 ( .A(n476), .B(n477), .ZN(SUM[11]) );
  NAND2_X1 U236 ( .A1(n472), .A2(n478), .ZN(n477) );
  NAND2_X1 U237 ( .A1(n473), .A2(n469), .ZN(n476) );
  NAND2_X1 U238 ( .A1(n475), .A2(n479), .ZN(n478) );
  XNOR2_X1 U239 ( .A(n80), .B(n81), .ZN(SUM[8]) );
  NAND2_X1 U240 ( .A1(n82), .A2(n83), .ZN(n80) );
  XNOR2_X1 U241 ( .A(n467), .B(n466), .ZN(SUM[12]) );
  NAND2_X1 U242 ( .A1(n449), .A2(n440), .ZN(n467) );
  XNOR2_X1 U243 ( .A(n421), .B(n575), .ZN(SUM[1]) );
  NAND2_X1 U244 ( .A1(n352), .A2(n351), .ZN(n421) );
  XNOR2_X1 U245 ( .A(n123), .B(n97), .ZN(SUM[5]) );
  NAND2_X1 U246 ( .A1(n96), .A2(n95), .ZN(n123) );
  XNOR2_X1 U247 ( .A(n92), .B(n90), .ZN(SUM[6]) );
  NAND2_X1 U248 ( .A1(n91), .A2(n88), .ZN(n92) );
  XNOR2_X1 U249 ( .A(n76), .B(n77), .ZN(SUM[9]) );
  NAND2_X1 U250 ( .A1(n78), .A2(n79), .ZN(n76) );
  XNOR2_X1 U251 ( .A(n480), .B(n479), .ZN(SUM[10]) );
  NAND2_X1 U252 ( .A1(n475), .A2(n472), .ZN(n480) );
  XNOR2_X1 U253 ( .A(n349), .B(n284), .ZN(SUM[2]) );
  NAND2_X1 U254 ( .A1(n285), .A2(n282), .ZN(n349) );
  XNOR2_X1 U255 ( .A(n201), .B(n455), .ZN(SUM[4]) );
  NAND2_X1 U256 ( .A1(n126), .A2(n125), .ZN(n201) );
  OAI21_X1 U257 ( .B1(n490), .B2(n491), .A(n281), .ZN(n455) );
  NAND2_X1 U258 ( .A1(n285), .A2(n280), .ZN(n491) );
  NOR2_X1 U259 ( .A1(n492), .A2(n493), .ZN(n490) );
  NAND2_X1 U260 ( .A1(n282), .A2(n351), .ZN(n493) );
  OAI21_X1 U261 ( .B1(n567), .B2(n566), .A(n79), .ZN(n479) );
  INV_X1 U262 ( .A(n77), .ZN(n567) );
  INV_X1 U263 ( .A(n78), .ZN(n566) );
  OAI21_X1 U264 ( .B1(n563), .B2(n562), .A(n441), .ZN(n460) );
  INV_X1 U265 ( .A(n463), .ZN(n563) );
  OAI21_X1 U266 ( .B1(n400), .B2(n553), .A(n391), .ZN(n398) );
  OAI21_X1 U267 ( .B1(n571), .B2(n573), .A(n125), .ZN(n97) );
  INV_X1 U268 ( .A(n126), .ZN(n571) );
  OAI21_X1 U269 ( .B1(n549), .B2(n551), .A(n368), .ZN(n377) );
  INV_X1 U270 ( .A(n369), .ZN(n549) );
  OAI21_X1 U271 ( .B1(n570), .B2(n569), .A(n95), .ZN(n90) );
  INV_X1 U272 ( .A(n96), .ZN(n569) );
  INV_X1 U273 ( .A(n97), .ZN(n570) );
  OAI21_X1 U274 ( .B1(n548), .B2(n547), .A(n367), .ZN(n373) );
  INV_X1 U275 ( .A(n364), .ZN(n547) );
  INV_X1 U276 ( .A(n377), .ZN(n548) );
  OAI21_X1 U277 ( .B1(n559), .B2(n558), .A(n415), .ZN(n426) );
  INV_X1 U278 ( .A(n429), .ZN(n559) );
  NAND4_X1 U279 ( .A1(n393), .A2(n389), .A3(n390), .A4(n385), .ZN(n335) );
  NAND4_X1 U280 ( .A1(n369), .A2(n364), .A3(n366), .A4(n361), .ZN(n329) );
  OAI21_X1 U281 ( .B1(n407), .B2(n408), .A(n409), .ZN(n332) );
  NAND2_X1 U282 ( .A1(n410), .A2(n411), .ZN(n408) );
  NOR2_X1 U283 ( .A1(n412), .A2(n413), .ZN(n407) );
  NAND2_X1 U284 ( .A1(n414), .A2(n415), .ZN(n413) );
  OAI21_X1 U285 ( .B1(n383), .B2(n384), .A(n385), .ZN(n334) );
  NAND2_X1 U286 ( .A1(n386), .A2(n387), .ZN(n384) );
  NOR2_X1 U287 ( .A1(n16), .A2(n388), .ZN(n383) );
  AND2_X1 U288 ( .A1(n391), .A2(n392), .ZN(n16) );
  OAI21_X1 U289 ( .B1(n15), .B2(n360), .A(n361), .ZN(n330) );
  AND3_X1 U290 ( .A1(n364), .A2(n365), .A3(n366), .ZN(n15) );
  NAND2_X1 U291 ( .A1(n362), .A2(n363), .ZN(n360) );
  NAND2_X1 U292 ( .A1(n367), .A2(n368), .ZN(n365) );
  NAND4_X1 U293 ( .A1(n418), .A2(n419), .A3(n410), .A4(n411), .ZN(n341) );
  NAND4_X1 U294 ( .A1(n126), .A2(n96), .A3(n91), .A4(n86), .ZN(n456) );
  NAND4_X1 U295 ( .A1(n78), .A2(n82), .A3(n475), .A4(n469), .ZN(n454) );
  OAI211_X1 U296 ( .C1(n562), .C2(n440), .A(n441), .B(n442), .ZN(n436) );
  NOR2_X1 U297 ( .A1(n558), .A2(n417), .ZN(n412) );
  NOR2_X1 U298 ( .A1(n574), .A2(n422), .ZN(n492) );
  INV_X1 U299 ( .A(n352), .ZN(n574) );
  NAND2_X1 U300 ( .A1(n483), .A2(n83), .ZN(n77) );
  NAND2_X1 U301 ( .A1(n81), .A2(n82), .ZN(n483) );
  NAND2_X1 U302 ( .A1(n465), .A2(n440), .ZN(n463) );
  NAND2_X1 U303 ( .A1(n466), .A2(n449), .ZN(n465) );
  NAND2_X1 U304 ( .A1(n431), .A2(n417), .ZN(n429) );
  NAND2_X1 U305 ( .A1(n420), .A2(n418), .ZN(n431) );
  NAND2_X1 U306 ( .A1(n350), .A2(n351), .ZN(n284) );
  NAND2_X1 U307 ( .A1(n352), .A2(n575), .ZN(n350) );
  OAI21_X1 U308 ( .B1(n514), .B2(n535), .A(net431068), .ZN(net431064) );
  INV_X1 U309 ( .A(net431069), .ZN(n535) );
  INV_X1 U310 ( .A(net538409), .ZN(n514) );
  NAND2_X1 U311 ( .A1(n469), .A2(n470), .ZN(n451) );
  NAND2_X1 U312 ( .A1(n79), .A2(n83), .ZN(n474) );
  NAND2_X1 U313 ( .A1(n86), .A2(n484), .ZN(n453) );
  NAND2_X1 U314 ( .A1(n95), .A2(n125), .ZN(n486) );
  INV_X1 U315 ( .A(n422), .ZN(n575) );
  AND2_X1 U316 ( .A1(n404), .A2(n392), .ZN(n400) );
  NAND2_X1 U317 ( .A1(n394), .A2(n393), .ZN(n404) );
  AND4_X1 U318 ( .A1(n339), .A2(n340), .A3(n325), .A4(n326), .ZN(n72) );
  INV_X1 U319 ( .A(n419), .ZN(n558) );
  INV_X1 U320 ( .A(n450), .ZN(n562) );
  NAND2_X1 U321 ( .A1(n389), .A2(n390), .ZN(n388) );
  AND4_X1 U322 ( .A1(n449), .A2(n450), .A3(n443), .A4(n444), .ZN(n14) );
  AND2_X1 U323 ( .A1(n444), .A2(n443), .ZN(n435) );
  INV_X1 U324 ( .A(n438), .ZN(n561) );
  NAND2_X1 U325 ( .A1(A[52]), .A2(B[52]), .ZN(n158) );
  NOR2_X1 U326 ( .A1(A[53]), .A2(B[53]), .ZN(n157) );
  NAND2_X1 U327 ( .A1(n149), .A2(n12), .ZN(n193) );
  XOR2_X1 U328 ( .A(n127), .B(n129), .Z(SUM[59]) );
  OR2_X1 U329 ( .A1(A[34]), .A2(B[34]), .ZN(n298) );
  NOR2_X1 U330 ( .A1(A[29]), .A2(B[29]), .ZN(n3) );
  OAI21_X1 U331 ( .B1(n266), .B2(n521), .A(n267), .ZN(n224) );
  INV_X1 U332 ( .A(n270), .ZN(n521) );
  OAI211_X1 U333 ( .C1(A[38]), .C2(B[38]), .A(n271), .B(n272), .ZN(n270) );
  NOR2_X1 U334 ( .A1(B[49]), .A2(A[49]), .ZN(n188) );
  NAND2_X1 U335 ( .A1(B[45]), .A2(A[45]), .ZN(n212) );
  NAND2_X1 U336 ( .A1(B[41]), .A2(A[41]), .ZN(n251) );
  NAND2_X1 U337 ( .A1(B[52]), .A2(A[52]), .ZN(n168) );
  NAND2_X1 U338 ( .A1(B[36]), .A2(A[36]), .ZN(n275) );
  NAND2_X1 U339 ( .A1(B[40]), .A2(A[40]), .ZN(n252) );
  OR2_X1 U340 ( .A1(A[35]), .A2(B[35]), .ZN(n299) );
  NAND2_X1 U341 ( .A1(B[32]), .A2(A[32]), .ZN(n305) );
  NAND2_X1 U342 ( .A1(A[38]), .A2(B[38]), .ZN(n269) );
  OR2_X1 U343 ( .A1(B[37]), .A2(A[37]), .ZN(n271) );
  OR2_X1 U344 ( .A1(B[33]), .A2(A[33]), .ZN(n297) );
  OAI21_X1 U345 ( .B1(n33), .B2(n209), .A(n210), .ZN(n207) );
  AOI21_X1 U346 ( .B1(n211), .B2(n212), .A(n56), .ZN(n209) );
  NOR2_X1 U347 ( .A1(B[46]), .A2(A[46]), .ZN(n56) );
  NAND2_X1 U348 ( .A1(n526), .A2(n215), .ZN(n211) );
  OR2_X1 U349 ( .A1(B[32]), .A2(A[32]), .ZN(n296) );
  NAND2_X1 U350 ( .A1(B[29]), .A2(A[29]), .ZN(n323) );
  OR2_X1 U351 ( .A1(B[30]), .A2(A[30]), .ZN(n325) );
  OR2_X1 U352 ( .A1(B[26]), .A2(A[26]), .ZN(n366) );
  NAND2_X1 U353 ( .A1(B[34]), .A2(A[34]), .ZN(n307) );
  NAND2_X1 U354 ( .A1(B[33]), .A2(A[33]), .ZN(n306) );
  OAI21_X1 U355 ( .B1(B[59]), .B2(A[59]), .A(n112), .ZN(n111) );
  OR2_X1 U356 ( .A1(B[25]), .A2(A[25]), .ZN(n364) );
  NAND2_X1 U357 ( .A1(B[30]), .A2(A[30]), .ZN(n324) );
  NAND2_X1 U358 ( .A1(B[37]), .A2(A[37]), .ZN(n274) );
  NAND2_X1 U359 ( .A1(B[49]), .A2(A[49]), .ZN(n190) );
  NAND2_X1 U360 ( .A1(A[58]), .A2(B[58]), .ZN(n119) );
  OR2_X1 U361 ( .A1(A[31]), .A2(B[31]), .ZN(n326) );
  NAND2_X1 U362 ( .A1(B[42]), .A2(A[42]), .ZN(n246) );
  NAND2_X1 U363 ( .A1(B[56]), .A2(A[56]), .ZN(n139) );
  NAND2_X1 U364 ( .A1(B[28]), .A2(A[28]), .ZN(n322) );
  OR2_X1 U365 ( .A1(B[36]), .A2(A[36]), .ZN(n276) );
  NAND2_X1 U366 ( .A1(A[48]), .A2(B[48]), .ZN(n189) );
  OR2_X1 U367 ( .A1(B[41]), .A2(A[41]), .ZN(n248) );
  OR2_X1 U368 ( .A1(B[27]), .A2(A[27]), .ZN(n361) );
  NAND2_X1 U369 ( .A1(A[59]), .A2(B[59]), .ZN(n118) );
  OR2_X1 U370 ( .A1(A[58]), .A2(B[58]), .ZN(n112) );
  NAND2_X1 U371 ( .A1(B[44]), .A2(A[44]), .ZN(n216) );
  OR2_X1 U372 ( .A1(B[28]), .A2(A[28]), .ZN(n339) );
  OR2_X1 U373 ( .A1(B[21]), .A2(A[21]), .ZN(n389) );
  OR2_X1 U374 ( .A1(B[56]), .A2(A[56]), .ZN(n113) );
  NAND2_X1 U375 ( .A1(A[50]), .A2(B[50]), .ZN(n191) );
  OR2_X1 U376 ( .A1(A[38]), .A2(B[38]), .ZN(n273) );
  OR2_X1 U377 ( .A1(A[46]), .A2(B[46]), .ZN(n213) );
  NAND2_X1 U378 ( .A1(B[31]), .A2(A[31]), .ZN(n320) );
  OR2_X1 U379 ( .A1(A[47]), .A2(B[47]), .ZN(n210) );
  OR2_X1 U380 ( .A1(B[44]), .A2(A[44]), .ZN(n227) );
  NAND2_X1 U381 ( .A1(B[35]), .A2(A[35]), .ZN(n302) );
  OR2_X1 U382 ( .A1(B[39]), .A2(A[39]), .ZN(n267) );
  AND2_X1 U383 ( .A1(A[46]), .A2(B[46]), .ZN(n33) );
  OR2_X1 U384 ( .A1(A[48]), .A2(B[48]), .ZN(n185) );
  OR2_X1 U385 ( .A1(B[40]), .A2(A[40]), .ZN(n254) );
  OR2_X1 U386 ( .A1(A[29]), .A2(B[29]), .ZN(n340) );
  OR2_X1 U387 ( .A1(A[43]), .A2(B[43]), .ZN(n243) );
  NAND2_X1 U388 ( .A1(n114), .A2(n74), .ZN(n120) );
  AND2_X1 U389 ( .A1(A[56]), .A2(B[56]), .ZN(n74) );
  OR2_X1 U390 ( .A1(B[22]), .A2(A[22]), .ZN(n390) );
  OR2_X1 U391 ( .A1(B[18]), .A2(A[18]), .ZN(n410) );
  OR2_X1 U392 ( .A1(B[14]), .A2(A[14]), .ZN(n443) );
  OR2_X1 U393 ( .A1(B[19]), .A2(A[19]), .ZN(n411) );
  OR2_X1 U394 ( .A1(B[23]), .A2(A[23]), .ZN(n385) );
  OR2_X1 U395 ( .A1(B[16]), .A2(A[16]), .ZN(n418) );
  OR2_X1 U396 ( .A1(B[17]), .A2(A[17]), .ZN(n419) );
  OR2_X1 U397 ( .A1(B[13]), .A2(A[13]), .ZN(n450) );
  OR2_X1 U398 ( .A1(B[20]), .A2(A[20]), .ZN(n393) );
  OR2_X1 U399 ( .A1(B[24]), .A2(A[24]), .ZN(n369) );
  OR2_X1 U400 ( .A1(B[15]), .A2(A[15]), .ZN(n444) );
  OR2_X1 U401 ( .A1(B[6]), .A2(A[6]), .ZN(n91) );
  OR2_X1 U402 ( .A1(B[10]), .A2(A[10]), .ZN(n475) );
  OR2_X1 U403 ( .A1(B[5]), .A2(A[5]), .ZN(n96) );
  OR2_X1 U404 ( .A1(B[9]), .A2(A[9]), .ZN(n78) );
  OR2_X1 U405 ( .A1(B[11]), .A2(A[11]), .ZN(n469) );
  OR2_X1 U406 ( .A1(B[7]), .A2(A[7]), .ZN(n86) );
  OR2_X1 U407 ( .A1(B[8]), .A2(A[8]), .ZN(n82) );
  OR2_X1 U408 ( .A1(B[2]), .A2(A[2]), .ZN(n285) );
  OR2_X1 U409 ( .A1(B[12]), .A2(A[12]), .ZN(n449) );
  OR2_X1 U410 ( .A1(B[1]), .A2(A[1]), .ZN(n352) );
  OR2_X1 U411 ( .A1(B[4]), .A2(A[4]), .ZN(n126) );
  OR2_X1 U412 ( .A1(B[3]), .A2(A[3]), .ZN(n280) );
  OR2_X1 U413 ( .A1(B[0]), .A2(A[0]), .ZN(n489) );
  INV_X1 U414 ( .A(B[54]), .ZN(n572) );
  NAND2_X1 U415 ( .A1(B[8]), .A2(A[8]), .ZN(n83) );
  NAND2_X1 U416 ( .A1(B[1]), .A2(A[1]), .ZN(n351) );
  NAND2_X1 U417 ( .A1(B[12]), .A2(A[12]), .ZN(n440) );
  NAND2_X1 U418 ( .A1(B[14]), .A2(A[14]), .ZN(n442) );
  NAND2_X1 U419 ( .A1(B[4]), .A2(A[4]), .ZN(n125) );
  NAND2_X1 U420 ( .A1(B[24]), .A2(A[24]), .ZN(n368) );
  NAND2_X1 U421 ( .A1(B[17]), .A2(A[17]), .ZN(n415) );
  NAND2_X1 U422 ( .A1(B[13]), .A2(A[13]), .ZN(n441) );
  NAND2_X1 U423 ( .A1(B[26]), .A2(A[26]), .ZN(n363) );
  NAND2_X1 U424 ( .A1(B[22]), .A2(A[22]), .ZN(n387) );
  NAND2_X1 U425 ( .A1(B[16]), .A2(A[16]), .ZN(n417) );
  NAND2_X1 U426 ( .A1(B[5]), .A2(A[5]), .ZN(n95) );
  NAND2_X1 U427 ( .A1(B[9]), .A2(A[9]), .ZN(n79) );
  NAND2_X1 U428 ( .A1(B[25]), .A2(A[25]), .ZN(n367) );
  NAND2_X1 U429 ( .A1(B[18]), .A2(A[18]), .ZN(n414) );
  NAND2_X1 U430 ( .A1(B[2]), .A2(A[2]), .ZN(n282) );
  NAND2_X1 U431 ( .A1(B[0]), .A2(A[0]), .ZN(n422) );
  NAND2_X1 U432 ( .A1(B[6]), .A2(A[6]), .ZN(n88) );
  NAND2_X1 U433 ( .A1(B[10]), .A2(A[10]), .ZN(n472) );
  NAND2_X1 U434 ( .A1(B[21]), .A2(A[21]), .ZN(n391) );
  NAND2_X1 U435 ( .A1(B[20]), .A2(A[20]), .ZN(n392) );
  NAND2_X1 U436 ( .A1(B[3]), .A2(A[3]), .ZN(n281) );
  NAND2_X1 U437 ( .A1(B[27]), .A2(A[27]), .ZN(n362) );
  NAND2_X1 U438 ( .A1(B[15]), .A2(A[15]), .ZN(n438) );
  NAND2_X1 U439 ( .A1(B[19]), .A2(A[19]), .ZN(n409) );
  NAND2_X1 U440 ( .A1(B[23]), .A2(A[23]), .ZN(n386) );
  NAND2_X1 U441 ( .A1(B[7]), .A2(A[7]), .ZN(n87) );
  NAND2_X1 U442 ( .A1(B[11]), .A2(A[11]), .ZN(n473) );
  OR2_X1 U443 ( .A1(A[55]), .A2(B[55]), .ZN(n156) );
  XNOR2_X1 U444 ( .A(n178), .B(n177), .ZN(SUM[53]) );
  NAND2_X1 U445 ( .A1(n179), .A2(n168), .ZN(n178) );
  XNOR2_X1 U446 ( .A(n194), .B(n193), .ZN(SUM[51]) );
  NAND2_X1 U447 ( .A1(n195), .A2(n191), .ZN(n194) );
  NAND2_X1 U448 ( .A1(B[51]), .A2(n503), .ZN(n149) );
  NOR2_X1 U449 ( .A1(A[51]), .A2(B[51]), .ZN(n68) );
  OR2_X1 U450 ( .A1(n503), .A2(B[51]), .ZN(n12) );
  NAND2_X1 U451 ( .A1(n242), .A2(n220), .ZN(n240) );
  OAI21_X1 U452 ( .B1(n219), .B2(n525), .A(n220), .ZN(n218) );
  AND2_X1 U453 ( .A1(n220), .A2(n216), .ZN(n65) );
  NAND2_X1 U454 ( .A1(n143), .A2(n109), .ZN(n141) );
  NOR2_X1 U455 ( .A1(n151), .A2(n152), .ZN(n146) );
  OR2_X1 U456 ( .A1(A[59]), .A2(B[59]), .ZN(n62) );
  AND2_X1 U457 ( .A1(B[60]), .A2(A[60]), .ZN(net537977) );
  NAND2_X1 U458 ( .A1(B[60]), .A2(A[60]), .ZN(net431068) );
  NOR2_X1 U459 ( .A1(n134), .A2(n541), .ZN(n130) );
  XNOR2_X1 U460 ( .A(n28), .B(n204), .ZN(SUM[48]) );
  NAND2_X1 U461 ( .A1(n40), .A2(n147), .ZN(n42) );
  NOR2_X1 U462 ( .A1(n151), .A2(n152), .ZN(n40) );
  NAND2_X1 U463 ( .A1(n155), .A2(n156), .ZN(n151) );
  AND2_X1 U464 ( .A1(n62), .A2(n112), .ZN(n115) );
  NAND2_X1 U465 ( .A1(n120), .A2(n71), .ZN(n116) );
  XNOR2_X1 U466 ( .A(n499), .B(n263), .ZN(SUM[40]) );
  NAND2_X1 U467 ( .A1(n253), .A2(n21), .ZN(n242) );
  NAND2_X1 U468 ( .A1(n253), .A2(n254), .ZN(n262) );
  NOR2_X1 U469 ( .A1(n111), .A2(n134), .ZN(n104) );
  INV_X1 U470 ( .A(n115), .ZN(n530) );
  AOI21_X1 U471 ( .B1(n115), .B2(n116), .A(n531), .ZN(n102) );
  NAND2_X1 U472 ( .A1(n185), .A2(n189), .ZN(n204) );
  NAND2_X1 U473 ( .A1(n197), .A2(n189), .ZN(n203) );
  INV_X1 U474 ( .A(n189), .ZN(n528) );
  OAI211_X1 U475 ( .C1(n188), .C2(n189), .A(n190), .B(n191), .ZN(n187) );
  OR2_X1 U476 ( .A1(B[63]), .A2(A[63]), .ZN(n100) );
  INV_X1 U477 ( .A(n39), .ZN(n534) );
  OR2_X1 U478 ( .A1(B[62]), .A2(A[62]), .ZN(n39) );
  INV_X1 U479 ( .A(n165), .ZN(n512) );
  NAND2_X1 U480 ( .A1(n63), .A2(n64), .ZN(n58) );
  NAND2_X1 U481 ( .A1(n242), .A2(n65), .ZN(n63) );
  XNOR2_X1 U482 ( .A(n233), .B(n232), .ZN(SUM[47]) );
  NAND2_X1 U483 ( .A1(n234), .A2(n524), .ZN(n233) );
  XNOR2_X1 U484 ( .A(n144), .B(n131), .ZN(SUM[56]) );
  AOI21_X1 U485 ( .B1(n130), .B2(n131), .A(n132), .ZN(n127) );
  NAND2_X1 U486 ( .A1(n46), .A2(n185), .ZN(n197) );
  XNOR2_X1 U487 ( .A(n287), .B(n286), .ZN(SUM[39]) );
  XNOR2_X1 U488 ( .A(n289), .B(n290), .ZN(SUM[38]) );
  NAND2_X1 U489 ( .A1(n273), .A2(n289), .ZN(n288) );
  INV_X1 U490 ( .A(n110), .ZN(n538) );
  AOI21_X1 U491 ( .B1(n60), .B2(n110), .A(n30), .ZN(n145) );
  AOI21_X1 U492 ( .B1(n60), .B2(n110), .A(n30), .ZN(n143) );
  INV_X1 U493 ( .A(n231), .ZN(n522) );
  XNOR2_X1 U494 ( .A(n135), .B(n136), .ZN(SUM[58]) );
  NAND2_X1 U495 ( .A1(n42), .A2(n145), .ZN(n131) );
  OAI211_X1 U496 ( .C1(n157), .C2(n158), .A(n159), .B(n160), .ZN(n110) );
  NAND2_X1 U497 ( .A1(A[53]), .A2(B[53]), .ZN(n159) );
  AOI21_X1 U498 ( .B1(n141), .B2(n113), .A(n532), .ZN(n140) );
  NAND2_X1 U499 ( .A1(n235), .A2(n213), .ZN(n234) );
  NAND2_X1 U500 ( .A1(n247), .A2(n243), .ZN(n255) );
  NAND2_X1 U501 ( .A1(n243), .A2(n244), .ZN(n220) );
  NAND2_X1 U502 ( .A1(A[43]), .A2(B[43]), .ZN(n247) );
  NAND2_X1 U503 ( .A1(n533), .A2(n35), .ZN(n36) );
  NAND2_X1 U504 ( .A1(n114), .A2(n113), .ZN(n134) );
  XNOR2_X1 U505 ( .A(n36), .B(net431081), .ZN(SUM[62]) );
  NAND2_X1 U506 ( .A1(net431064), .A2(net431065), .ZN(net431061) );
  OR2_X1 U507 ( .A1(A[61]), .A2(B[61]), .ZN(net431065) );
  NAND2_X1 U508 ( .A1(net431059), .A2(n38), .ZN(net431057) );
  NAND2_X1 U509 ( .A1(n39), .A2(n38), .ZN(net431081) );
  XNOR2_X1 U510 ( .A(n140), .B(n8), .ZN(SUM[57]) );
  XNOR2_X1 U511 ( .A(n166), .B(n180), .ZN(SUM[52]) );
  AOI21_X1 U512 ( .B1(n166), .B2(n153), .A(n167), .ZN(n165) );
  NAND2_X1 U513 ( .A1(n166), .A2(n153), .ZN(n179) );
  NAND2_X1 U514 ( .A1(n186), .A2(n187), .ZN(n148) );
  AND2_X1 U515 ( .A1(n114), .A2(n121), .ZN(n8) );
  OAI21_X1 U516 ( .B1(n138), .B2(n139), .A(n121), .ZN(n47) );
  OAI211_X1 U517 ( .C1(n1), .C2(n530), .A(n103), .B(n118), .ZN(net538409) );
  OAI21_X1 U518 ( .B1(n498), .B2(B[59]), .A(n118), .ZN(n129) );
  INV_X1 U519 ( .A(n118), .ZN(n531) );
  NAND2_X1 U521 ( .A1(n537), .A2(n572), .ZN(n161) );
  NAND2_X1 U522 ( .A1(n537), .A2(n572), .ZN(n154) );
  NAND2_X1 U523 ( .A1(n268), .A2(n267), .ZN(n286) );
  NAND2_X1 U524 ( .A1(n268), .A2(n269), .ZN(n266) );
  NAND2_X1 U525 ( .A1(n104), .A2(n105), .ZN(n103) );
  AND2_X1 U526 ( .A1(A[55]), .A2(B[55]), .ZN(n30) );
  OR2_X1 U527 ( .A1(B[55]), .A2(A[55]), .ZN(n66) );
  INV_X1 U528 ( .A(n150), .ZN(n511) );
  NAND2_X1 U529 ( .A1(n181), .A2(n150), .ZN(n166) );
  NAND4_X1 U530 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n46) );
  NAND4_X1 U531 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n28) );
  AOI21_X1 U532 ( .B1(net431070), .B2(net431069), .A(net537977), .ZN(net431086) );
  XNOR2_X1 U533 ( .A(net431072), .B(n101), .ZN(SUM[63]) );
  OAI21_X1 U536 ( .B1(net431073), .B2(n534), .A(n38), .ZN(net431072) );
  AOI21_X1 U537 ( .B1(n131), .B2(n61), .A(n496), .ZN(n135) );
  NAND2_X1 U538 ( .A1(n47), .A2(n112), .ZN(n133) );
  NOR2_X1 U539 ( .A1(B[57]), .A2(A[57]), .ZN(n138) );
  NAND2_X1 U540 ( .A1(A[57]), .A2(B[57]), .ZN(n121) );
  XNOR2_X1 U541 ( .A(net431086), .B(net431087), .ZN(SUM[61]) );
  NAND2_X1 U542 ( .A1(B[47]), .A2(n497), .ZN(n208) );
  OR2_X1 U543 ( .A1(A[47]), .A2(B[47]), .ZN(n226) );
  OAI21_X1 U544 ( .B1(n99), .B2(net431057), .A(n100), .ZN(n98) );
  NAND2_X1 U545 ( .A1(net431059), .A2(n100), .ZN(n101) );
  XNOR2_X1 U546 ( .A(n504), .B(n196), .ZN(SUM[50]) );
  NAND2_X1 U547 ( .A1(n24), .A2(n543), .ZN(n195) );
  NAND2_X1 U548 ( .A1(A[62]), .A2(B[62]), .ZN(n38) );
  AOI21_X1 U549 ( .B1(net431061), .B2(n34), .A(n534), .ZN(n99) );
  AND2_X1 U550 ( .A1(n34), .A2(net431065), .ZN(net431087) );
  OAI21_X1 U551 ( .B1(net431068), .B2(n37), .A(n34), .ZN(net431076) );
  NOR2_X1 U552 ( .A1(n57), .A2(n505), .ZN(n183) );
  NOR2_X1 U553 ( .A1(n68), .A2(n57), .ZN(n186) );
  AND2_X1 U554 ( .A1(B[54]), .A2(A[54]), .ZN(n73) );
  NAND2_X1 U555 ( .A1(A[54]), .A2(B[54]), .ZN(n160) );
  INV_X1 U556 ( .A(A[54]), .ZN(n537) );
  NAND2_X1 U557 ( .A1(n23), .A2(n250), .ZN(n257) );
  INV_X1 U558 ( .A(n224), .ZN(n520) );
  NAND2_X1 U559 ( .A1(A[39]), .A2(B[39]), .ZN(n268) );
  NOR2_X1 U560 ( .A1(n515), .A2(net431076), .ZN(net431073) );
  INV_X1 U561 ( .A(net431076), .ZN(n533) );
  NAND2_X1 U562 ( .A1(A[61]), .A2(B[61]), .ZN(n34) );
  NOR2_X1 U563 ( .A1(B[61]), .A2(A[61]), .ZN(n37) );
  NAND2_X1 U564 ( .A1(n146), .A2(n147), .ZN(n109) );
  NAND2_X1 U565 ( .A1(n102), .A2(n103), .ZN(net431070) );
  NAND2_X1 U566 ( .A1(B[63]), .A2(A[63]), .ZN(net431059) );
endmodule


module RCA_NBIT64_2 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_2_DW01_add_3 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module RCA_NBIT64_1_DW01_add_4 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   net430041, net430036, net430025, net430023, net430018, net430017,
         net430011, net430005, net430003, net430001, net429999, net429979,
         net429975, net429974, net429968, net534717, net534765, net537145,
         net430016, net537152, net535584, net429988, net429987, net429982,
         net429972, net429970, net429969, net429989, net429973, net429991,
         net429990, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14,
         n16, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n34,
         n37, n38, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51, n52, n55,
         n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n101,
         n102, n104, n105, n106, n107, n108, n109, n112, n113, n114, n117,
         n118, n119, n120, n122, n123, n124, n125, n126, n127, n128, n129,
         n133, n134, n135, n136, n137, n138, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n151, n153, n155, n156, n157, n158,
         n160, n161, n162, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n179, n180, n181, n182, n184,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n219,
         n220, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n247, n248, n249, n250, n251, n252, n253, n254,
         n256, n257, n258, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n289, n291, n292,
         n293, n296, n297, n298, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n311, n313, n314, n315, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n334, n335, n337, n338, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n359, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n386, n387, n388, n389, n390, n391, n392, n393, n395, n397,
         n398, n399, n400, n401, n404, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n440, n441, n442, n443, n446, n447, n448, n449,
         n450, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526;

  NAND3_X1 U51 ( .A1(n129), .A2(n472), .A3(n128), .ZN(n37) );
  NAND3_X1 U485 ( .A1(n95), .A2(n94), .A3(n93), .ZN(net430003) );
  NAND3_X1 U496 ( .A1(n129), .A2(n472), .A3(n128), .ZN(n95) );
  NAND3_X1 U502 ( .A1(n149), .A2(n148), .A3(n147), .ZN(n146) );
  NAND3_X1 U547 ( .A1(n428), .A2(n429), .A3(n430), .ZN(n427) );
  NAND3_X1 U548 ( .A1(n431), .A2(n67), .A3(n432), .ZN(n428) );
  NAND3_X1 U553 ( .A1(n442), .A2(n77), .A3(n76), .ZN(n441) );
  NAND3_X1 U554 ( .A1(n85), .A2(n443), .A3(n80), .ZN(n442) );
  OR2_X1 U2 ( .A1(A[59]), .A2(B[59]), .ZN(net430036) );
  AND2_X1 U3 ( .A1(n446), .A2(n379), .ZN(SUM[0]) );
  CLKBUF_X1 U4 ( .A(A[47]), .Z(n453) );
  CLKBUF_X1 U5 ( .A(A[59]), .Z(n454) );
  OAI21_X1 U6 ( .B1(n8), .B2(n204), .A(n205), .ZN(n455) );
  CLKBUF_X1 U7 ( .A(n92), .Z(n456) );
  BUF_X1 U8 ( .A(net535584), .Z(n457) );
  NOR2_X1 U9 ( .A1(A[61]), .A2(B[61]), .ZN(net535584) );
  CLKBUF_X1 U10 ( .A(A[57]), .Z(n458) );
  AND2_X1 U11 ( .A1(n166), .A2(n151), .ZN(n459) );
  AND2_X1 U12 ( .A1(n160), .A2(n459), .ZN(n149) );
  OR2_X2 U13 ( .A1(B[42]), .A2(A[42]), .ZN(n210) );
  XNOR2_X1 U14 ( .A(net429982), .B(n460), .ZN(SUM[63]) );
  AND2_X1 U15 ( .A1(net429972), .A2(n47), .ZN(n460) );
  XOR2_X1 U16 ( .A(n19), .B(n461), .Z(SUM[41]) );
  NAND2_X1 U17 ( .A1(n208), .A2(n211), .ZN(n461) );
  INV_X1 U18 ( .A(n232), .ZN(n469) );
  INV_X1 U19 ( .A(n337), .ZN(n502) );
  INV_X1 U20 ( .A(n377), .ZN(n511) );
  NAND2_X1 U21 ( .A1(n28), .A2(n213), .ZN(n203) );
  OR2_X1 U22 ( .A1(n188), .A2(n61), .ZN(n232) );
  AND2_X1 U23 ( .A1(n62), .A2(n193), .ZN(n61) );
  AND2_X1 U24 ( .A1(n146), .A2(n145), .ZN(n143) );
  INV_X1 U25 ( .A(A[58]), .ZN(n477) );
  INV_X1 U26 ( .A(n117), .ZN(n476) );
  OAI21_X1 U27 ( .B1(n524), .B2(n413), .A(n410), .ZN(n70) );
  OAI21_X1 U28 ( .B1(n511), .B2(n298), .A(n507), .ZN(n351) );
  INV_X1 U29 ( .A(n289), .ZN(n507) );
  OAI21_X1 U30 ( .B1(n506), .B2(n292), .A(n291), .ZN(n337) );
  INV_X1 U31 ( .A(n351), .ZN(n506) );
  OAI21_X1 U32 ( .B1(n502), .B2(n286), .A(n287), .ZN(n314) );
  NAND4_X1 U33 ( .A1(n293), .A2(n508), .A3(n497), .A4(n63), .ZN(n272) );
  INV_X1 U34 ( .A(n298), .ZN(n508) );
  INV_X1 U35 ( .A(n286), .ZN(n497) );
  NOR2_X1 U36 ( .A1(n511), .A2(n292), .ZN(n293) );
  AOI21_X1 U37 ( .B1(n409), .B2(n410), .A(n411), .ZN(n404) );
  NAND2_X1 U38 ( .A1(n519), .A2(n412), .ZN(n409) );
  INV_X1 U39 ( .A(n413), .ZN(n519) );
  NAND2_X1 U40 ( .A1(n390), .A2(n391), .ZN(n377) );
  OAI21_X1 U41 ( .B1(n404), .B2(n516), .A(n10), .ZN(n390) );
  AOI21_X1 U42 ( .B1(n392), .B2(n393), .A(n512), .ZN(n391) );
  INV_X1 U43 ( .A(n408), .ZN(n516) );
  NAND2_X1 U44 ( .A1(n425), .A2(n408), .ZN(n423) );
  NAND2_X1 U45 ( .A1(n515), .A2(n70), .ZN(n425) );
  INV_X1 U46 ( .A(n411), .ZN(n515) );
  NAND2_X1 U47 ( .A1(n63), .A2(n284), .ZN(n273) );
  OAI21_X1 U48 ( .B1(n285), .B2(n286), .A(n287), .ZN(n284) );
  AOI21_X1 U49 ( .B1(n501), .B2(n289), .A(n503), .ZN(n285) );
  INV_X1 U50 ( .A(n291), .ZN(n503) );
  INV_X1 U52 ( .A(n412), .ZN(n524) );
  INV_X1 U53 ( .A(n292), .ZN(n501) );
  INV_X1 U54 ( .A(net429968), .ZN(SUM[64]) );
  OAI21_X1 U55 ( .B1(n13), .B2(n471), .A(n261), .ZN(n266) );
  AND2_X1 U56 ( .A1(n270), .A2(n260), .ZN(n13) );
  OAI21_X1 U57 ( .B1(n16), .B2(n494), .A(n229), .ZN(n244) );
  AND2_X1 U58 ( .A1(n249), .A2(n230), .ZN(n16) );
  INV_X1 U59 ( .A(n226), .ZN(n494) );
  AND3_X1 U60 ( .A1(n208), .A2(n209), .A3(n210), .ZN(n8) );
  NAND2_X1 U61 ( .A1(n211), .A2(n212), .ZN(n209) );
  OAI21_X1 U62 ( .B1(n25), .B2(n493), .A(n180), .ZN(n196) );
  AND2_X1 U63 ( .A1(n200), .A2(n179), .ZN(n25) );
  AOI21_X1 U64 ( .B1(n91), .B2(n57), .A(net534765), .ZN(n89) );
  INV_X1 U65 ( .A(n64), .ZN(n473) );
  OAI21_X1 U66 ( .B1(n222), .B2(n7), .A(n1), .ZN(n189) );
  AND3_X1 U67 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n7) );
  NAND2_X1 U68 ( .A1(n224), .A2(n225), .ZN(n222) );
  NAND2_X1 U69 ( .A1(n229), .A2(n230), .ZN(n227) );
  OAI21_X1 U70 ( .B1(n470), .B2(n256), .A(n257), .ZN(n188) );
  INV_X1 U71 ( .A(n258), .ZN(n470) );
  NAND2_X1 U72 ( .A1(n254), .A2(n253), .ZN(n256) );
  OAI211_X1 U73 ( .C1(n471), .C2(n260), .A(n261), .B(n262), .ZN(n258) );
  AOI21_X1 U74 ( .B1(n122), .B2(n97), .A(n481), .ZN(n124) );
  AOI21_X1 U75 ( .B1(n153), .B2(n488), .A(n489), .ZN(n145) );
  INV_X1 U76 ( .A(n155), .ZN(n489) );
  OAI211_X1 U77 ( .C1(n491), .C2(n156), .A(n157), .B(n158), .ZN(n153) );
  INV_X1 U78 ( .A(n43), .ZN(n488) );
  AOI21_X1 U79 ( .B1(n57), .B2(n91), .A(net534765), .ZN(n92) );
  NAND4_X1 U80 ( .A1(n272), .A2(n273), .A3(n274), .A4(n275), .ZN(n14) );
  AND2_X1 U81 ( .A1(n29), .A2(n14), .ZN(n190) );
  AND4_X1 U82 ( .A1(n1), .A2(n226), .A3(n228), .A4(n231), .ZN(n29) );
  OAI21_X1 U83 ( .B1(n30), .B2(n491), .A(n157), .ZN(n164) );
  AND2_X1 U84 ( .A1(n170), .A2(n156), .ZN(n30) );
  INV_X1 U85 ( .A(n188), .ZN(n468) );
  OAI21_X1 U86 ( .B1(n143), .B2(n474), .A(n134), .ZN(n56) );
  OAI21_X1 U87 ( .B1(n19), .B2(n492), .A(n211), .ZN(n22) );
  NAND4_X1 U88 ( .A1(n272), .A2(n273), .A3(n274), .A4(n275), .ZN(n193) );
  AOI21_X1 U89 ( .B1(net430023), .B2(net430016), .A(n484), .ZN(net430017) );
  AOI21_X1 U90 ( .B1(n109), .B2(n108), .A(n479), .ZN(n106) );
  INV_X1 U91 ( .A(net429999), .ZN(n479) );
  NOR2_X1 U92 ( .A1(n476), .A2(n487), .ZN(n108) );
  OAI21_X1 U93 ( .B1(n59), .B2(n480), .A(n112), .ZN(n109) );
  AND2_X1 U94 ( .A1(n93), .A2(n94), .ZN(n127) );
  AND2_X1 U95 ( .A1(n219), .A2(n212), .ZN(n19) );
  NAND2_X1 U96 ( .A1(n2), .A2(n214), .ZN(n219) );
  NAND2_X1 U97 ( .A1(net430036), .A2(net430041), .ZN(n51) );
  NOR2_X1 U98 ( .A1(net534717), .A2(net430001), .ZN(n50) );
  OAI21_X1 U99 ( .B1(n464), .B2(n490), .A(n158), .ZN(n162) );
  INV_X1 U100 ( .A(n147), .ZN(n490) );
  INV_X1 U101 ( .A(n97), .ZN(n480) );
  INV_X1 U102 ( .A(n98), .ZN(n487) );
  NOR2_X1 U103 ( .A1(n487), .A2(n480), .ZN(n123) );
  INV_X1 U104 ( .A(n297), .ZN(n495) );
  AND3_X1 U105 ( .A1(n37), .A2(n94), .A3(n93), .ZN(n59) );
  XNOR2_X1 U106 ( .A(n119), .B(n118), .ZN(SUM[58]) );
  NAND2_X1 U107 ( .A1(n117), .A2(net429999), .ZN(n118) );
  NOR2_X1 U108 ( .A1(net534765), .A2(n482), .ZN(n107) );
  NAND2_X1 U109 ( .A1(n276), .A2(n277), .ZN(n274) );
  OAI211_X1 U110 ( .C1(n495), .C2(n279), .A(n280), .B(n281), .ZN(n277) );
  AND2_X1 U111 ( .A1(n283), .A2(n282), .ZN(n276) );
  INV_X1 U112 ( .A(n144), .ZN(n474) );
  INV_X1 U113 ( .A(n114), .ZN(n481) );
  AND2_X1 U114 ( .A1(net430036), .A2(net430041), .ZN(n57) );
  INV_X1 U115 ( .A(n140), .ZN(n475) );
  NAND2_X1 U116 ( .A1(n193), .A2(n251), .ZN(n270) );
  NAND2_X1 U117 ( .A1(n232), .A2(n231), .ZN(n249) );
  OAI21_X1 U118 ( .B1(n143), .B2(n474), .A(n134), .ZN(n141) );
  NAND2_X1 U119 ( .A1(n201), .A2(n191), .ZN(n200) );
  NAND2_X1 U120 ( .A1(n270), .A2(n260), .ZN(n268) );
  NAND2_X1 U121 ( .A1(n155), .A2(n160), .ZN(n161) );
  XNOR2_X1 U122 ( .A(n27), .B(n26), .ZN(SUM[47]) );
  AND2_X1 U123 ( .A1(n175), .A2(n23), .ZN(n26) );
  XNOR2_X1 U124 ( .A(n56), .B(n142), .ZN(SUM[53]) );
  NAND2_X1 U125 ( .A1(n140), .A2(n135), .ZN(n142) );
  NAND2_X1 U126 ( .A1(n147), .A2(n158), .ZN(n165) );
  XNOR2_X1 U127 ( .A(n143), .B(n24), .ZN(SUM[52]) );
  AND2_X1 U128 ( .A1(n134), .A2(n144), .ZN(n24) );
  XNOR2_X1 U129 ( .A(n196), .B(n197), .ZN(SUM[46]) );
  NAND2_X1 U130 ( .A1(n182), .A2(n181), .ZN(n197) );
  XNOR2_X1 U131 ( .A(n167), .B(n169), .ZN(SUM[49]) );
  NAND2_X1 U132 ( .A1(n166), .A2(n157), .ZN(n169) );
  XNOR2_X1 U133 ( .A(n21), .B(n20), .ZN(SUM[43]) );
  XNOR2_X1 U134 ( .A(n198), .B(n199), .ZN(SUM[45]) );
  NAND2_X1 U135 ( .A1(n192), .A2(n180), .ZN(n199) );
  NAND2_X1 U136 ( .A1(n156), .A2(n151), .ZN(n171) );
  XNOR2_X1 U137 ( .A(n22), .B(n217), .ZN(SUM[42]) );
  NAND2_X1 U138 ( .A1(n210), .A2(n207), .ZN(n217) );
  XNOR2_X1 U139 ( .A(n201), .B(n202), .ZN(SUM[44]) );
  NAND2_X1 U140 ( .A1(n191), .A2(n179), .ZN(n202) );
  XNOR2_X1 U141 ( .A(n213), .B(n220), .ZN(SUM[40]) );
  NAND2_X1 U142 ( .A1(n214), .A2(n212), .ZN(n220) );
  XNOR2_X1 U143 ( .A(n267), .B(n266), .ZN(SUM[34]) );
  NAND2_X1 U144 ( .A1(n253), .A2(n262), .ZN(n267) );
  XNOR2_X1 U145 ( .A(n263), .B(n264), .ZN(SUM[35]) );
  NAND2_X1 U146 ( .A1(n257), .A2(n254), .ZN(n264) );
  XNOR2_X1 U147 ( .A(n242), .B(n241), .ZN(SUM[39]) );
  NAND2_X1 U148 ( .A1(n224), .A2(n1), .ZN(n241) );
  XNOR2_X1 U149 ( .A(n244), .B(n245), .ZN(SUM[38]) );
  NAND2_X1 U150 ( .A1(n228), .A2(n225), .ZN(n245) );
  XNOR2_X1 U151 ( .A(n248), .B(n247), .ZN(SUM[37]) );
  NAND2_X1 U152 ( .A1(n249), .A2(n230), .ZN(n247) );
  XNOR2_X1 U153 ( .A(n250), .B(n232), .ZN(SUM[36]) );
  NAND2_X1 U154 ( .A1(n231), .A2(n230), .ZN(n250) );
  XNOR2_X1 U155 ( .A(n357), .B(n359), .ZN(SUM[21]) );
  NOR2_X1 U156 ( .A1(n505), .A2(n504), .ZN(n359) );
  XNOR2_X1 U157 ( .A(n335), .B(n334), .ZN(SUM[25]) );
  NAND2_X1 U158 ( .A1(n321), .A2(n324), .ZN(n335) );
  XNOR2_X1 U159 ( .A(n331), .B(n330), .ZN(SUM[26]) );
  NAND2_X1 U160 ( .A1(n323), .A2(n320), .ZN(n331) );
  XNOR2_X1 U161 ( .A(n327), .B(n328), .ZN(SUM[27]) );
  NAND2_X1 U162 ( .A1(n320), .A2(n329), .ZN(n327) );
  XNOR2_X1 U163 ( .A(n315), .B(n314), .ZN(SUM[28]) );
  NAND2_X1 U164 ( .A1(n296), .A2(n279), .ZN(n315) );
  XNOR2_X1 U165 ( .A(n305), .B(n311), .ZN(SUM[29]) );
  NOR2_X1 U166 ( .A1(n496), .A2(n495), .ZN(n311) );
  XNOR2_X1 U167 ( .A(n304), .B(n303), .ZN(SUM[30]) );
  NAND2_X1 U168 ( .A1(n282), .A2(n281), .ZN(n304) );
  XNOR2_X1 U169 ( .A(n300), .B(n301), .ZN(SUM[31]) );
  NAND2_X1 U170 ( .A1(n281), .A2(n302), .ZN(n301) );
  XNOR2_X1 U171 ( .A(n269), .B(n268), .ZN(SUM[33]) );
  NAND2_X1 U172 ( .A1(n252), .A2(n261), .ZN(n269) );
  NOR2_X1 U173 ( .A1(n486), .A2(net537152), .ZN(net430005) );
  XNOR2_X1 U174 ( .A(n55), .B(net430025), .ZN(SUM[60]) );
  NAND2_X1 U175 ( .A1(net430016), .A2(net430011), .ZN(net430025) );
  AND2_X1 U176 ( .A1(n94), .A2(n137), .ZN(n38) );
  XNOR2_X1 U177 ( .A(n124), .B(n125), .ZN(SUM[57]) );
  NOR2_X1 U178 ( .A1(net534717), .A2(n487), .ZN(n125) );
  XNOR2_X1 U179 ( .A(n4), .B(n34), .ZN(SUM[54]) );
  OR2_X1 U180 ( .A1(n64), .A2(n6), .ZN(n34) );
  XNOR2_X1 U181 ( .A(n59), .B(n126), .ZN(SUM[56]) );
  NOR2_X1 U182 ( .A1(n481), .A2(n480), .ZN(n126) );
  XNOR2_X1 U183 ( .A(n271), .B(n14), .ZN(SUM[32]) );
  NAND2_X1 U184 ( .A1(n260), .A2(n251), .ZN(n271) );
  INV_X1 U185 ( .A(n346), .ZN(n504) );
  INV_X1 U186 ( .A(n208), .ZN(n492) );
  INV_X1 U187 ( .A(net430011), .ZN(n484) );
  INV_X1 U188 ( .A(n252), .ZN(n471) );
  NAND2_X1 U189 ( .A1(n170), .A2(n156), .ZN(n167) );
  INV_X1 U190 ( .A(n166), .ZN(n491) );
  INV_X1 U191 ( .A(n192), .ZN(n493) );
  NAND2_X1 U192 ( .A1(n200), .A2(n179), .ZN(n198) );
  NAND2_X1 U193 ( .A1(n243), .A2(n225), .ZN(n242) );
  NAND2_X1 U194 ( .A1(n228), .A2(n244), .ZN(n243) );
  NAND2_X1 U195 ( .A1(n226), .A2(n229), .ZN(n248) );
  NAND2_X1 U196 ( .A1(n275), .A2(n283), .ZN(n300) );
  NAND2_X1 U197 ( .A1(n262), .A2(n265), .ZN(n263) );
  NAND2_X1 U198 ( .A1(n266), .A2(n253), .ZN(n265) );
  NAND2_X1 U199 ( .A1(n176), .A2(n177), .ZN(n174) );
  OAI211_X1 U200 ( .C1(n493), .C2(n179), .A(n180), .B(n181), .ZN(n177) );
  AND2_X1 U201 ( .A1(n23), .A2(n182), .ZN(n176) );
  NAND2_X1 U202 ( .A1(n318), .A2(n319), .ZN(n328) );
  INV_X1 U203 ( .A(net429973), .ZN(n486) );
  NAND2_X1 U204 ( .A1(n3), .A2(n184), .ZN(n173) );
  AND4_X1 U205 ( .A1(n254), .A2(n252), .A3(n253), .A4(n251), .ZN(n62) );
  AND2_X1 U206 ( .A1(n195), .A2(n181), .ZN(n27) );
  NAND2_X1 U207 ( .A1(n196), .A2(n182), .ZN(n195) );
  AND2_X1 U208 ( .A1(n215), .A2(n207), .ZN(n21) );
  NAND2_X1 U209 ( .A1(n210), .A2(n216), .ZN(n215) );
  OAI21_X1 U210 ( .B1(n19), .B2(n492), .A(n211), .ZN(n216) );
  INV_X1 U211 ( .A(net429975), .ZN(n485) );
  AND2_X1 U212 ( .A1(n98), .A2(n60), .ZN(net430001) );
  AND2_X1 U213 ( .A1(n113), .A2(n114), .ZN(n112) );
  INV_X1 U214 ( .A(net430016), .ZN(n483) );
  INV_X1 U215 ( .A(net430036), .ZN(n482) );
  INV_X1 U216 ( .A(net537145), .ZN(n478) );
  XNOR2_X1 U217 ( .A(n421), .B(n420), .ZN(SUM[13]) );
  NAND2_X1 U218 ( .A1(n407), .A2(n398), .ZN(n421) );
  XNOR2_X1 U219 ( .A(n414), .B(n415), .ZN(SUM[15]) );
  NAND2_X1 U220 ( .A1(n416), .A2(n399), .ZN(n415) );
  XNOR2_X1 U221 ( .A(n389), .B(n377), .ZN(SUM[16]) );
  NAND2_X1 U222 ( .A1(n374), .A2(n375), .ZN(n389) );
  XNOR2_X1 U223 ( .A(n387), .B(n386), .ZN(SUM[17]) );
  NAND2_X1 U224 ( .A1(n376), .A2(n372), .ZN(n387) );
  XNOR2_X1 U225 ( .A(n384), .B(n383), .ZN(SUM[18]) );
  NAND2_X1 U226 ( .A1(n367), .A2(n371), .ZN(n384) );
  XNOR2_X1 U227 ( .A(n380), .B(n381), .ZN(SUM[19]) );
  NAND2_X1 U228 ( .A1(n371), .A2(n382), .ZN(n380) );
  XNOR2_X1 U229 ( .A(n362), .B(n351), .ZN(SUM[20]) );
  NAND2_X1 U230 ( .A1(n350), .A2(n349), .ZN(n362) );
  XNOR2_X1 U231 ( .A(n356), .B(n355), .ZN(SUM[22]) );
  NAND2_X1 U232 ( .A1(n347), .A2(n344), .ZN(n356) );
  XNOR2_X1 U233 ( .A(n352), .B(n353), .ZN(SUM[23]) );
  NAND2_X1 U234 ( .A1(n344), .A2(n354), .ZN(n353) );
  XNOR2_X1 U235 ( .A(n338), .B(n337), .ZN(SUM[24]) );
  NAND2_X1 U236 ( .A1(n326), .A2(n325), .ZN(n338) );
  NAND2_X1 U237 ( .A1(n366), .A2(n368), .ZN(n381) );
  NAND2_X1 U238 ( .A1(n343), .A2(n342), .ZN(n352) );
  NAND2_X1 U239 ( .A1(n395), .A2(n401), .ZN(n414) );
  XNOR2_X1 U240 ( .A(n418), .B(n417), .ZN(SUM[14]) );
  NAND2_X1 U241 ( .A1(n400), .A2(n399), .ZN(n418) );
  XNOR2_X1 U242 ( .A(n69), .B(n70), .ZN(SUM[8]) );
  NAND2_X1 U243 ( .A1(n71), .A2(n72), .ZN(n69) );
  XNOR2_X1 U244 ( .A(n437), .B(n436), .ZN(SUM[10]) );
  NAND2_X1 U245 ( .A1(n432), .A2(n429), .ZN(n437) );
  XNOR2_X1 U246 ( .A(n233), .B(n234), .ZN(SUM[3]) );
  NAND2_X1 U247 ( .A1(n237), .A2(n238), .ZN(n233) );
  NAND2_X1 U248 ( .A1(n235), .A2(n236), .ZN(n234) );
  NAND2_X1 U249 ( .A1(n239), .A2(n240), .ZN(n238) );
  XNOR2_X1 U250 ( .A(n306), .B(n239), .ZN(SUM[2]) );
  NAND2_X1 U251 ( .A1(n240), .A2(n237), .ZN(n306) );
  XNOR2_X1 U252 ( .A(n81), .B(n79), .ZN(SUM[6]) );
  NAND2_X1 U253 ( .A1(n80), .A2(n77), .ZN(n81) );
  XNOR2_X1 U254 ( .A(n73), .B(n74), .ZN(SUM[7]) );
  NAND2_X1 U255 ( .A1(n77), .A2(n78), .ZN(n73) );
  XNOR2_X1 U256 ( .A(n65), .B(n66), .ZN(SUM[9]) );
  NAND2_X1 U257 ( .A1(n67), .A2(n68), .ZN(n65) );
  XNOR2_X1 U258 ( .A(n433), .B(n434), .ZN(SUM[11]) );
  NAND2_X1 U259 ( .A1(n429), .A2(n435), .ZN(n434) );
  XNOR2_X1 U260 ( .A(n424), .B(n423), .ZN(SUM[12]) );
  NAND2_X1 U261 ( .A1(n406), .A2(n397), .ZN(n424) );
  XNOR2_X1 U262 ( .A(n378), .B(n526), .ZN(SUM[1]) );
  NAND2_X1 U263 ( .A1(n309), .A2(n308), .ZN(n378) );
  XNOR2_X1 U264 ( .A(n168), .B(n412), .ZN(SUM[4]) );
  NAND2_X1 U265 ( .A1(n105), .A2(n104), .ZN(n168) );
  XNOR2_X1 U266 ( .A(n102), .B(n86), .ZN(SUM[5]) );
  NAND2_X1 U267 ( .A1(n85), .A2(n84), .ZN(n102) );
  NAND2_X1 U268 ( .A1(n430), .A2(n426), .ZN(n433) );
  NAND2_X1 U269 ( .A1(n75), .A2(n76), .ZN(n74) );
  OAI21_X1 U270 ( .B1(n447), .B2(n448), .A(n236), .ZN(n412) );
  NAND2_X1 U271 ( .A1(n240), .A2(n235), .ZN(n448) );
  NOR2_X1 U272 ( .A1(n449), .A2(n450), .ZN(n447) );
  NAND2_X1 U273 ( .A1(n237), .A2(n308), .ZN(n450) );
  OAI21_X1 U274 ( .B1(n518), .B2(n517), .A(n68), .ZN(n436) );
  INV_X1 U275 ( .A(n66), .ZN(n518) );
  INV_X1 U276 ( .A(n67), .ZN(n517) );
  OAI21_X1 U277 ( .B1(n514), .B2(n513), .A(n398), .ZN(n417) );
  INV_X1 U278 ( .A(n420), .ZN(n514) );
  OAI21_X1 U279 ( .B1(n357), .B2(n504), .A(n348), .ZN(n355) );
  OAI21_X1 U280 ( .B1(n305), .B2(n495), .A(n280), .ZN(n303) );
  OAI21_X1 U281 ( .B1(n522), .B2(n524), .A(n104), .ZN(n86) );
  INV_X1 U282 ( .A(n105), .ZN(n522) );
  OAI21_X1 U283 ( .B1(n500), .B2(n502), .A(n325), .ZN(n334) );
  INV_X1 U284 ( .A(n326), .ZN(n500) );
  OAI21_X1 U285 ( .B1(n521), .B2(n520), .A(n84), .ZN(n79) );
  INV_X1 U286 ( .A(n85), .ZN(n520) );
  INV_X1 U287 ( .A(n86), .ZN(n521) );
  OAI21_X1 U288 ( .B1(n510), .B2(n509), .A(n372), .ZN(n383) );
  INV_X1 U289 ( .A(n386), .ZN(n510) );
  OAI21_X1 U290 ( .B1(n499), .B2(n498), .A(n324), .ZN(n330) );
  INV_X1 U291 ( .A(n321), .ZN(n498) );
  INV_X1 U292 ( .A(n334), .ZN(n499) );
  NAND4_X1 U293 ( .A1(n347), .A2(n350), .A3(n342), .A4(n346), .ZN(n292) );
  NAND4_X1 U294 ( .A1(n326), .A2(n321), .A3(n323), .A4(n318), .ZN(n286) );
  OAI21_X1 U295 ( .B1(n364), .B2(n365), .A(n366), .ZN(n289) );
  NAND2_X1 U296 ( .A1(n367), .A2(n368), .ZN(n365) );
  NOR2_X1 U297 ( .A1(n369), .A2(n370), .ZN(n364) );
  NAND2_X1 U298 ( .A1(n371), .A2(n372), .ZN(n370) );
  NAND2_X1 U299 ( .A1(net429972), .A2(net429973), .ZN(net429970) );
  AOI21_X1 U300 ( .B1(net429974), .B2(net429975), .A(net537152), .ZN(net429969) );
  OAI21_X1 U301 ( .B1(n484), .B2(n55), .A(net429979), .ZN(net429974) );
  OAI21_X1 U302 ( .B1(n340), .B2(n341), .A(n342), .ZN(n291) );
  NAND2_X1 U303 ( .A1(n343), .A2(n344), .ZN(n341) );
  NOR2_X1 U304 ( .A1(n12), .A2(n345), .ZN(n340) );
  AND2_X1 U305 ( .A1(n348), .A2(n349), .ZN(n12) );
  OAI21_X1 U306 ( .B1(n11), .B2(n317), .A(n318), .ZN(n287) );
  AND3_X1 U307 ( .A1(n321), .A2(n322), .A3(n323), .ZN(n11) );
  NAND2_X1 U308 ( .A1(n319), .A2(n320), .ZN(n317) );
  NAND2_X1 U309 ( .A1(n324), .A2(n325), .ZN(n322) );
  NAND4_X1 U310 ( .A1(n375), .A2(n376), .A3(n367), .A4(n368), .ZN(n298) );
  NAND4_X1 U311 ( .A1(n105), .A2(n85), .A3(n80), .A4(n75), .ZN(n413) );
  NAND4_X1 U312 ( .A1(n67), .A2(n71), .A3(n432), .A4(n426), .ZN(n411) );
  OAI211_X1 U313 ( .C1(n513), .C2(n397), .A(n398), .B(n399), .ZN(n393) );
  NOR2_X1 U314 ( .A1(n509), .A2(n374), .ZN(n369) );
  NOR2_X1 U315 ( .A1(n525), .A2(n379), .ZN(n449) );
  INV_X1 U316 ( .A(n309), .ZN(n525) );
  NAND2_X1 U317 ( .A1(n440), .A2(n72), .ZN(n66) );
  NAND2_X1 U318 ( .A1(n70), .A2(n71), .ZN(n440) );
  NAND2_X1 U319 ( .A1(n422), .A2(n397), .ZN(n420) );
  NAND2_X1 U320 ( .A1(n423), .A2(n406), .ZN(n422) );
  NAND2_X1 U321 ( .A1(n388), .A2(n374), .ZN(n386) );
  NAND2_X1 U322 ( .A1(n377), .A2(n375), .ZN(n388) );
  NAND2_X1 U323 ( .A1(n307), .A2(n308), .ZN(n239) );
  NAND2_X1 U324 ( .A1(n309), .A2(n526), .ZN(n307) );
  NAND2_X1 U325 ( .A1(n426), .A2(n427), .ZN(n408) );
  NAND2_X1 U326 ( .A1(n68), .A2(n72), .ZN(n431) );
  NAND2_X1 U327 ( .A1(n75), .A2(n441), .ZN(n410) );
  NAND2_X1 U328 ( .A1(n84), .A2(n104), .ZN(n443) );
  INV_X1 U329 ( .A(n379), .ZN(n526) );
  AND2_X1 U330 ( .A1(n313), .A2(n279), .ZN(n305) );
  NAND2_X1 U331 ( .A1(n314), .A2(n296), .ZN(n313) );
  AND2_X1 U332 ( .A1(n361), .A2(n349), .ZN(n357) );
  NAND2_X1 U333 ( .A1(n351), .A2(n350), .ZN(n361) );
  AND4_X1 U334 ( .A1(n296), .A2(n297), .A3(n282), .A4(n283), .ZN(n63) );
  NAND2_X1 U335 ( .A1(n79), .A2(n80), .ZN(n78) );
  NAND2_X1 U336 ( .A1(n383), .A2(n367), .ZN(n382) );
  NAND2_X1 U337 ( .A1(n330), .A2(n323), .ZN(n329) );
  INV_X1 U338 ( .A(n376), .ZN(n509) );
  INV_X1 U339 ( .A(n407), .ZN(n513) );
  NAND2_X1 U340 ( .A1(n282), .A2(n303), .ZN(n302) );
  NAND2_X1 U341 ( .A1(n347), .A2(n355), .ZN(n354) );
  NAND2_X1 U342 ( .A1(n432), .A2(n436), .ZN(n435) );
  NAND2_X1 U343 ( .A1(n346), .A2(n347), .ZN(n345) );
  NAND2_X1 U344 ( .A1(n400), .A2(n417), .ZN(n416) );
  AND4_X1 U345 ( .A1(n406), .A2(n407), .A3(n400), .A4(n401), .ZN(n10) );
  AND2_X1 U346 ( .A1(n401), .A2(n400), .ZN(n392) );
  INV_X1 U347 ( .A(n280), .ZN(n496) );
  INV_X1 U348 ( .A(n348), .ZN(n505) );
  INV_X1 U349 ( .A(n395), .ZN(n512) );
  NAND2_X1 U350 ( .A1(B[54]), .A2(A[54]), .ZN(n136) );
  NOR2_X1 U351 ( .A1(B[62]), .A2(A[62]), .ZN(net537152) );
  OR2_X1 U352 ( .A1(B[38]), .A2(A[38]), .ZN(n228) );
  NOR2_X1 U353 ( .A1(B[54]), .A2(A[54]), .ZN(n64) );
  OR2_X1 U354 ( .A1(B[37]), .A2(A[37]), .ZN(n226) );
  NAND4_X1 U355 ( .A1(n223), .A2(n226), .A3(n231), .A4(n228), .ZN(n194) );
  OR2_X1 U356 ( .A1(B[39]), .A2(A[39]), .ZN(n223) );
  NAND2_X1 U357 ( .A1(B[36]), .A2(A[36]), .ZN(n230) );
  NAND2_X1 U358 ( .A1(B[44]), .A2(A[44]), .ZN(n179) );
  OR2_X1 U359 ( .A1(A[36]), .A2(B[36]), .ZN(n231) );
  NAND2_X1 U360 ( .A1(B[48]), .A2(A[48]), .ZN(n156) );
  NAND2_X1 U361 ( .A1(B[32]), .A2(A[32]), .ZN(n260) );
  OR2_X1 U362 ( .A1(A[34]), .A2(B[34]), .ZN(n253) );
  NAND2_X1 U363 ( .A1(B[41]), .A2(A[41]), .ZN(n211) );
  NAND2_X1 U364 ( .A1(B[58]), .A2(A[58]), .ZN(net429999) );
  NAND2_X1 U365 ( .A1(B[31]), .A2(A[31]), .ZN(n275) );
  AND2_X1 U366 ( .A1(n454), .A2(B[59]), .ZN(net534765) );
  NAND2_X1 U367 ( .A1(B[50]), .A2(A[50]), .ZN(n158) );
  NAND2_X1 U368 ( .A1(B[38]), .A2(A[38]), .ZN(n225) );
  OR2_X1 U369 ( .A1(B[26]), .A2(A[26]), .ZN(n323) );
  NAND2_X1 U370 ( .A1(B[52]), .A2(A[52]), .ZN(n134) );
  NAND2_X1 U371 ( .A1(B[49]), .A2(A[49]), .ZN(n157) );
  NAND2_X1 U372 ( .A1(B[33]), .A2(A[33]), .ZN(n261) );
  NAND2_X1 U373 ( .A1(B[45]), .A2(A[45]), .ZN(n180) );
  OR2_X1 U374 ( .A1(B[30]), .A2(A[30]), .ZN(n282) );
  OR2_X1 U375 ( .A1(B[25]), .A2(A[25]), .ZN(n321) );
  NAND2_X1 U376 ( .A1(B[34]), .A2(A[34]), .ZN(n262) );
  NAND2_X1 U377 ( .A1(B[30]), .A2(A[30]), .ZN(n281) );
  NAND2_X1 U378 ( .A1(B[37]), .A2(A[37]), .ZN(n229) );
  NAND2_X1 U379 ( .A1(A[60]), .A2(B[60]), .ZN(net430011) );
  NAND2_X1 U380 ( .A1(A[53]), .A2(B[53]), .ZN(n135) );
  OR2_X1 U381 ( .A1(A[57]), .A2(B[57]), .ZN(n98) );
  NAND2_X1 U382 ( .A1(B[40]), .A2(A[40]), .ZN(n212) );
  OR2_X1 U383 ( .A1(A[32]), .A2(B[32]), .ZN(n251) );
  OR2_X1 U384 ( .A1(A[46]), .A2(B[46]), .ZN(n182) );
  NAND2_X1 U385 ( .A1(B[46]), .A2(A[46]), .ZN(n181) );
  OR2_X1 U386 ( .A1(B[56]), .A2(A[56]), .ZN(n97) );
  OR2_X1 U387 ( .A1(B[41]), .A2(A[41]), .ZN(n208) );
  OR2_X1 U388 ( .A1(B[21]), .A2(A[21]), .ZN(n346) );
  OR2_X1 U389 ( .A1(B[27]), .A2(A[27]), .ZN(n318) );
  OR2_X1 U390 ( .A1(B[39]), .A2(A[39]), .ZN(n1) );
  OR2_X1 U391 ( .A1(A[60]), .A2(B[60]), .ZN(net430016) );
  OR2_X1 U392 ( .A1(B[40]), .A2(A[40]), .ZN(n214) );
  OR2_X1 U393 ( .A1(B[28]), .A2(A[28]), .ZN(n296) );
  OR2_X1 U394 ( .A1(A[33]), .A2(B[33]), .ZN(n252) );
  OR2_X1 U395 ( .A1(A[35]), .A2(B[35]), .ZN(n254) );
  NAND2_X1 U396 ( .A1(B[42]), .A2(A[42]), .ZN(n207) );
  OR2_X1 U397 ( .A1(A[31]), .A2(B[31]), .ZN(n283) );
  NAND2_X1 U398 ( .A1(A[35]), .A2(B[35]), .ZN(n257) );
  NAND2_X1 U399 ( .A1(B[39]), .A2(A[39]), .ZN(n224) );
  OR2_X1 U400 ( .A1(B[50]), .A2(A[50]), .ZN(n147) );
  OR2_X1 U401 ( .A1(B[44]), .A2(A[44]), .ZN(n191) );
  NAND2_X1 U402 ( .A1(B[47]), .A2(n453), .ZN(n175) );
  OR2_X1 U403 ( .A1(B[49]), .A2(A[49]), .ZN(n166) );
  OR2_X1 U404 ( .A1(B[45]), .A2(A[45]), .ZN(n192) );
  NAND2_X1 U405 ( .A1(B[56]), .A2(A[56]), .ZN(n114) );
  OR2_X1 U406 ( .A1(B[48]), .A2(A[48]), .ZN(n151) );
  OR2_X1 U407 ( .A1(B[29]), .A2(A[29]), .ZN(n297) );
  OR2_X1 U408 ( .A1(A[53]), .A2(B[53]), .ZN(n140) );
  OR2_X1 U409 ( .A1(A[43]), .A2(B[43]), .ZN(n205) );
  AND4_X1 U410 ( .A1(net430036), .A2(n97), .A3(n98), .A4(n96), .ZN(net537145)
         );
  OR2_X1 U411 ( .A1(B[58]), .A2(A[58]), .ZN(n96) );
  NOR2_X1 U412 ( .A1(n462), .A2(n463), .ZN(n3) );
  NOR2_X1 U413 ( .A1(A[47]), .A2(B[47]), .ZN(n462) );
  NAND3_X1 U414 ( .A1(n182), .A2(n192), .A3(n191), .ZN(n463) );
  OR2_X1 U415 ( .A1(B[52]), .A2(A[52]), .ZN(n144) );
  AND2_X1 U416 ( .A1(A[56]), .A2(B[56]), .ZN(n60) );
  AND2_X1 U417 ( .A1(B[54]), .A2(A[54]), .ZN(n6) );
  OR2_X1 U418 ( .A1(A[47]), .A2(B[47]), .ZN(n23) );
  OR2_X1 U419 ( .A1(B[18]), .A2(A[18]), .ZN(n367) );
  OR2_X1 U420 ( .A1(B[22]), .A2(A[22]), .ZN(n347) );
  OR2_X1 U421 ( .A1(B[14]), .A2(A[14]), .ZN(n400) );
  OR2_X1 U422 ( .A1(B[19]), .A2(A[19]), .ZN(n368) );
  OR2_X1 U423 ( .A1(B[23]), .A2(A[23]), .ZN(n342) );
  OR2_X1 U424 ( .A1(B[16]), .A2(A[16]), .ZN(n375) );
  OR2_X1 U425 ( .A1(B[20]), .A2(A[20]), .ZN(n350) );
  OR2_X1 U426 ( .A1(B[17]), .A2(A[17]), .ZN(n376) );
  OR2_X1 U427 ( .A1(B[13]), .A2(A[13]), .ZN(n407) );
  OR2_X1 U428 ( .A1(B[24]), .A2(A[24]), .ZN(n326) );
  OR2_X1 U429 ( .A1(B[15]), .A2(A[15]), .ZN(n401) );
  OR2_X1 U430 ( .A1(B[6]), .A2(A[6]), .ZN(n80) );
  OR2_X1 U431 ( .A1(B[10]), .A2(A[10]), .ZN(n432) );
  OR2_X1 U432 ( .A1(B[5]), .A2(A[5]), .ZN(n85) );
  OR2_X1 U433 ( .A1(B[9]), .A2(A[9]), .ZN(n67) );
  OR2_X1 U434 ( .A1(B[11]), .A2(A[11]), .ZN(n426) );
  OR2_X1 U435 ( .A1(B[7]), .A2(A[7]), .ZN(n75) );
  OR2_X1 U436 ( .A1(B[8]), .A2(A[8]), .ZN(n71) );
  OR2_X1 U437 ( .A1(B[2]), .A2(A[2]), .ZN(n240) );
  OR2_X1 U438 ( .A1(B[12]), .A2(A[12]), .ZN(n406) );
  OR2_X1 U439 ( .A1(B[1]), .A2(A[1]), .ZN(n309) );
  OR2_X1 U440 ( .A1(B[4]), .A2(A[4]), .ZN(n105) );
  OR2_X1 U441 ( .A1(B[3]), .A2(A[3]), .ZN(n235) );
  INV_X1 U442 ( .A(B[58]), .ZN(n523) );
  OR2_X1 U443 ( .A1(B[0]), .A2(A[0]), .ZN(n446) );
  NAND2_X1 U444 ( .A1(B[8]), .A2(A[8]), .ZN(n72) );
  NAND2_X1 U445 ( .A1(B[1]), .A2(A[1]), .ZN(n308) );
  NAND2_X1 U446 ( .A1(B[12]), .A2(A[12]), .ZN(n397) );
  NAND2_X1 U447 ( .A1(B[14]), .A2(A[14]), .ZN(n399) );
  NAND2_X1 U448 ( .A1(B[4]), .A2(A[4]), .ZN(n104) );
  NAND2_X1 U449 ( .A1(B[17]), .A2(A[17]), .ZN(n372) );
  NAND2_X1 U450 ( .A1(B[24]), .A2(A[24]), .ZN(n325) );
  NAND2_X1 U451 ( .A1(B[13]), .A2(A[13]), .ZN(n398) );
  NAND2_X1 U452 ( .A1(B[22]), .A2(A[22]), .ZN(n344) );
  NAND2_X1 U453 ( .A1(B[26]), .A2(A[26]), .ZN(n320) );
  NAND2_X1 U454 ( .A1(B[16]), .A2(A[16]), .ZN(n374) );
  NAND2_X1 U455 ( .A1(B[29]), .A2(A[29]), .ZN(n280) );
  NAND2_X1 U456 ( .A1(B[5]), .A2(A[5]), .ZN(n84) );
  NAND2_X1 U457 ( .A1(B[9]), .A2(A[9]), .ZN(n68) );
  NAND2_X1 U458 ( .A1(B[25]), .A2(A[25]), .ZN(n324) );
  NAND2_X1 U459 ( .A1(B[18]), .A2(A[18]), .ZN(n371) );
  NAND2_X1 U460 ( .A1(B[2]), .A2(A[2]), .ZN(n237) );
  NAND2_X1 U461 ( .A1(B[0]), .A2(A[0]), .ZN(n379) );
  NAND2_X1 U462 ( .A1(B[28]), .A2(A[28]), .ZN(n279) );
  NAND2_X1 U463 ( .A1(B[6]), .A2(A[6]), .ZN(n77) );
  NAND2_X1 U464 ( .A1(B[10]), .A2(A[10]), .ZN(n429) );
  NAND2_X1 U465 ( .A1(B[21]), .A2(A[21]), .ZN(n348) );
  NAND2_X1 U466 ( .A1(B[20]), .A2(A[20]), .ZN(n349) );
  NAND2_X1 U467 ( .A1(B[3]), .A2(A[3]), .ZN(n236) );
  NAND2_X1 U468 ( .A1(B[27]), .A2(A[27]), .ZN(n319) );
  NAND2_X1 U469 ( .A1(B[15]), .A2(A[15]), .ZN(n395) );
  NAND2_X1 U470 ( .A1(B[19]), .A2(A[19]), .ZN(n366) );
  NAND2_X1 U471 ( .A1(B[23]), .A2(A[23]), .ZN(n343) );
  NAND2_X1 U472 ( .A1(B[7]), .A2(A[7]), .ZN(n76) );
  NAND2_X1 U473 ( .A1(B[11]), .A2(A[11]), .ZN(n430) );
  NAND2_X1 U474 ( .A1(n120), .A2(n113), .ZN(n119) );
  NAND4_X1 U475 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n52) );
  NAND4_X1 U476 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n148) );
  NAND4_X1 U477 ( .A1(n3), .A2(n62), .A3(n190), .A4(n28), .ZN(n172) );
  XNOR2_X1 U478 ( .A(n162), .B(n161), .ZN(SUM[51]) );
  XNOR2_X1 U479 ( .A(n52), .B(n171), .ZN(SUM[48]) );
  XNOR2_X1 U480 ( .A(n164), .B(n165), .ZN(SUM[50]) );
  INV_X1 U481 ( .A(n164), .ZN(n464) );
  NAND2_X1 U482 ( .A1(n52), .A2(n151), .ZN(n170) );
  AOI21_X1 U483 ( .B1(n138), .B2(n473), .A(n6), .ZN(n45) );
  OAI21_X1 U484 ( .B1(n122), .B2(n481), .A(n123), .ZN(n120) );
  NAND2_X1 U486 ( .A1(n127), .A2(n37), .ZN(n122) );
  INV_X1 U487 ( .A(n41), .ZN(n472) );
  NAND2_X1 U488 ( .A1(n146), .A2(n145), .ZN(n129) );
  OAI21_X1 U489 ( .B1(n5), .B2(n478), .A(n89), .ZN(n88) );
  OAI21_X1 U490 ( .B1(n469), .B2(n194), .A(n189), .ZN(n2) );
  OAI21_X1 U491 ( .B1(n469), .B2(n194), .A(n189), .ZN(n213) );
  INV_X1 U492 ( .A(n40), .ZN(n467) );
  OAI21_X1 U493 ( .B1(n194), .B2(n468), .A(n189), .ZN(n40) );
  AOI21_X1 U494 ( .B1(n50), .B2(net429999), .A(n51), .ZN(n49) );
  NAND2_X1 U495 ( .A1(n523), .A2(n477), .ZN(n117) );
  NAND2_X1 U497 ( .A1(n477), .A2(n523), .ZN(net430041) );
  AND4_X1 U498 ( .A1(n205), .A2(n208), .A3(n210), .A4(n214), .ZN(n28) );
  OAI21_X1 U499 ( .B1(n8), .B2(n204), .A(n205), .ZN(n187) );
  NAND4_X1 U500 ( .A1(n214), .A2(n208), .A3(n210), .A4(n205), .ZN(n186) );
  NAND2_X1 U501 ( .A1(B[63]), .A2(A[63]), .ZN(net429972) );
  OAI21_X1 U503 ( .B1(n465), .B2(n475), .A(n135), .ZN(n4) );
  OAI21_X1 U504 ( .B1(n465), .B2(n475), .A(n135), .ZN(n138) );
  NOR2_X1 U505 ( .A1(n475), .A2(n474), .ZN(n128) );
  OAI211_X1 U506 ( .C1(n475), .C2(n134), .A(n135), .B(n136), .ZN(n133) );
  AND2_X1 U507 ( .A1(n206), .A2(n205), .ZN(n20) );
  INV_X1 U508 ( .A(n141), .ZN(n465) );
  NAND2_X1 U509 ( .A1(n206), .A2(n207), .ZN(n204) );
  NAND2_X1 U510 ( .A1(A[43]), .A2(B[43]), .ZN(n206) );
  NAND2_X1 U511 ( .A1(net430003), .A2(net537145), .ZN(n90) );
  AND3_X1 U512 ( .A1(n95), .A2(n94), .A3(n93), .ZN(n5) );
  NAND2_X1 U513 ( .A1(n133), .A2(n472), .ZN(n93) );
  XNOR2_X1 U514 ( .A(n45), .B(n38), .ZN(SUM[55]) );
  OR2_X1 U515 ( .A1(A[51]), .A2(B[51]), .ZN(n160) );
  NAND2_X1 U516 ( .A1(A[51]), .A2(B[51]), .ZN(n155) );
  OAI22_X1 U517 ( .A1(A[51]), .A2(B[51]), .B1(B[50]), .B2(A[50]), .ZN(n43) );
  NAND2_X1 U518 ( .A1(A[62]), .A2(B[62]), .ZN(net429973) );
  OR2_X1 U519 ( .A1(A[62]), .A2(B[62]), .ZN(n46) );
  OAI21_X1 U520 ( .B1(n5), .B2(n478), .A(n48), .ZN(net429988) );
  OR2_X1 U521 ( .A1(A[55]), .A2(B[55]), .ZN(n137) );
  NAND2_X1 U522 ( .A1(A[55]), .A2(B[55]), .ZN(n94) );
  OAI22_X1 U523 ( .A1(A[55]), .A2(B[55]), .B1(B[54]), .B2(A[54]), .ZN(n41) );
  NOR2_X1 U524 ( .A1(n49), .A2(net534765), .ZN(n48) );
  NAND2_X1 U525 ( .A1(n458), .A2(B[57]), .ZN(n113) );
  AOI22_X1 U526 ( .A1(n98), .A2(n60), .B1(B[57]), .B2(n458), .ZN(n101) );
  AND2_X1 U527 ( .A1(B[57]), .A2(n458), .ZN(net534717) );
  XNOR2_X1 U528 ( .A(n106), .B(n107), .ZN(SUM[59]) );
  NAND2_X1 U529 ( .A1(n203), .A2(n455), .ZN(n201) );
  OAI21_X1 U530 ( .B1(n467), .B2(n186), .A(n187), .ZN(n184) );
  XNOR2_X1 U531 ( .A(n87), .B(net430005), .ZN(SUM[62]) );
  OAI21_X1 U532 ( .B1(net429969), .B2(net429970), .A(n47), .ZN(net429968) );
  XNOR2_X1 U533 ( .A(net430017), .B(net430018), .ZN(SUM[61]) );
  NAND2_X1 U534 ( .A1(n90), .A2(n456), .ZN(n55) );
  NAND2_X1 U535 ( .A1(n90), .A2(n92), .ZN(net430023) );
  NAND2_X1 U536 ( .A1(n101), .A2(net429999), .ZN(n91) );
  OR2_X1 U537 ( .A1(A[63]), .A2(B[63]), .ZN(n47) );
  NOR2_X1 U538 ( .A1(n485), .A2(n457), .ZN(net430018) );
  AOI21_X1 U539 ( .B1(n88), .B2(net429979), .A(net429991), .ZN(n87) );
  NOR2_X1 U540 ( .A1(n457), .A2(n483), .ZN(net429979) );
  NAND2_X1 U541 ( .A1(net429991), .A2(n46), .ZN(net429990) );
  OAI21_X1 U542 ( .B1(net535584), .B2(net430011), .A(net429975), .ZN(net429991) );
  NAND2_X1 U543 ( .A1(A[61]), .A2(B[61]), .ZN(net429975) );
  AOI21_X1 U544 ( .B1(net429988), .B2(net429987), .A(net429989), .ZN(net429982) );
  NAND2_X1 U545 ( .A1(net429990), .A2(net429973), .ZN(net429989) );
  NOR3_X1 U546 ( .A1(net537152), .A2(n483), .A3(n457), .ZN(net429987) );
endmodule


module RCA_NBIT64_1 ( A, B, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  output Co;


  RCA_NBIT64_1_DW01_add_4 r48 ( .A({1'b0, A}), .B({1'b0, B}), .CI(1'b0), .SUM(
        {Co, S}) );
endmodule


module FD_64 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;


  SDFF_X1 Q_reg ( .D(D), .SI(1'b0), .SE(RESET), .CK(CLK), .Q(Q) );
endmodule


module FD_63 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_62 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_61 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;


  SDFF_X1 Q_reg ( .D(D), .SI(1'b0), .SE(RESET), .CK(CLK), .Q(Q) );
endmodule


module FD_60 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_59 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_58 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_57 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_56 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_55 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_54 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_53 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_52 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_51 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_50 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_49 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_48 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_47 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_46 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_45 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_44 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_43 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_42 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_41 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_40 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_39 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_38 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_37 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_36 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_35 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_34 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_33 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_32 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_31 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_30 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_29 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_28 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_27 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_26 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_25 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_24 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_23 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_22 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_21 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_20 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_19 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_18 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_17 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_16 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_15 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_14 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_13 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_12 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_11 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_10 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_9 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_8 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_7 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_6 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(D), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n3), .ZN(N3) );
endmodule


module FD_5 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_4 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_3 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n3), .A2(RESET), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_2 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n3), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n3) );
endmodule


module FD_1 ( D, CLK, RESET, Q );
  input D, CLK, RESET;
  output Q;
  wire   N3, n3;

  DFF_X1 Q_reg ( .D(N3), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(RESET), .ZN(n3) );
  AND2_X1 U4 ( .A1(D), .A2(n3), .ZN(N3) );
endmodule


module FD_GENERIC_NBIT64 ( D, CLK, RESET, Q );
  input [63:0] D;
  output [63:0] Q;
  input CLK, RESET;
  wire   n13, n14, n15, n16, n17, n18, n19, n20;

  FD_64 FD_i_0 ( .D(D[0]), .CLK(CLK), .RESET(n20), .Q(Q[0]) );
  FD_63 FD_i_1 ( .D(D[1]), .CLK(CLK), .RESET(n15), .Q(Q[1]) );
  FD_62 FD_i_2 ( .D(D[2]), .CLK(CLK), .RESET(n19), .Q(Q[2]) );
  FD_61 FD_i_3 ( .D(D[3]), .CLK(CLK), .RESET(n20), .Q(Q[3]) );
  FD_60 FD_i_4 ( .D(D[4]), .CLK(CLK), .RESET(n20), .Q(Q[4]) );
  FD_59 FD_i_5 ( .D(D[5]), .CLK(CLK), .RESET(n20), .Q(Q[5]) );
  FD_58 FD_i_6 ( .D(D[6]), .CLK(CLK), .RESET(n19), .Q(Q[6]) );
  FD_57 FD_i_7 ( .D(D[7]), .CLK(CLK), .RESET(n19), .Q(Q[7]) );
  FD_56 FD_i_8 ( .D(D[8]), .CLK(CLK), .RESET(n19), .Q(Q[8]) );
  FD_55 FD_i_9 ( .D(D[9]), .CLK(CLK), .RESET(n19), .Q(Q[9]) );
  FD_54 FD_i_10 ( .D(D[10]), .CLK(CLK), .RESET(n19), .Q(Q[10]) );
  FD_53 FD_i_11 ( .D(D[11]), .CLK(CLK), .RESET(n19), .Q(Q[11]) );
  FD_52 FD_i_12 ( .D(D[12]), .CLK(CLK), .RESET(n19), .Q(Q[12]) );
  FD_51 FD_i_13 ( .D(D[13]), .CLK(CLK), .RESET(n19), .Q(Q[13]) );
  FD_50 FD_i_14 ( .D(D[14]), .CLK(CLK), .RESET(n19), .Q(Q[14]) );
  FD_49 FD_i_15 ( .D(D[15]), .CLK(CLK), .RESET(n19), .Q(Q[15]) );
  FD_48 FD_i_16 ( .D(D[16]), .CLK(CLK), .RESET(n18), .Q(Q[16]) );
  FD_47 FD_i_17 ( .D(D[17]), .CLK(CLK), .RESET(n19), .Q(Q[17]) );
  FD_46 FD_i_18 ( .D(D[18]), .CLK(CLK), .RESET(n18), .Q(Q[18]) );
  FD_45 FD_i_19 ( .D(D[19]), .CLK(CLK), .RESET(n18), .Q(Q[19]) );
  FD_44 FD_i_20 ( .D(D[20]), .CLK(CLK), .RESET(n18), .Q(Q[20]) );
  FD_43 FD_i_21 ( .D(D[21]), .CLK(CLK), .RESET(n18), .Q(Q[21]) );
  FD_42 FD_i_22 ( .D(D[22]), .CLK(CLK), .RESET(n18), .Q(Q[22]) );
  FD_41 FD_i_23 ( .D(D[23]), .CLK(CLK), .RESET(n18), .Q(Q[23]) );
  FD_40 FD_i_24 ( .D(D[24]), .CLK(CLK), .RESET(n18), .Q(Q[24]) );
  FD_39 FD_i_25 ( .D(D[25]), .CLK(CLK), .RESET(n18), .Q(Q[25]) );
  FD_38 FD_i_26 ( .D(D[26]), .CLK(CLK), .RESET(n18), .Q(Q[26]) );
  FD_37 FD_i_27 ( .D(D[27]), .CLK(CLK), .RESET(n18), .Q(Q[27]) );
  FD_36 FD_i_28 ( .D(D[28]), .CLK(CLK), .RESET(n18), .Q(Q[28]) );
  FD_35 FD_i_29 ( .D(D[29]), .CLK(CLK), .RESET(n17), .Q(Q[29]) );
  FD_34 FD_i_30 ( .D(D[30]), .CLK(CLK), .RESET(n17), .Q(Q[30]) );
  FD_33 FD_i_31 ( .D(D[31]), .CLK(CLK), .RESET(n17), .Q(Q[31]) );
  FD_32 FD_i_32 ( .D(D[32]), .CLK(CLK), .RESET(n15), .Q(Q[32]) );
  FD_31 FD_i_33 ( .D(D[33]), .CLK(CLK), .RESET(n17), .Q(Q[33]) );
  FD_30 FD_i_34 ( .D(D[34]), .CLK(CLK), .RESET(n17), .Q(Q[34]) );
  FD_29 FD_i_35 ( .D(D[35]), .CLK(CLK), .RESET(n17), .Q(Q[35]) );
  FD_28 FD_i_36 ( .D(D[36]), .CLK(CLK), .RESET(n17), .Q(Q[36]) );
  FD_27 FD_i_37 ( .D(D[37]), .CLK(CLK), .RESET(n17), .Q(Q[37]) );
  FD_26 FD_i_38 ( .D(D[38]), .CLK(CLK), .RESET(n16), .Q(Q[38]) );
  FD_25 FD_i_39 ( .D(D[39]), .CLK(CLK), .RESET(n16), .Q(Q[39]) );
  FD_24 FD_i_40 ( .D(D[40]), .CLK(CLK), .RESET(n16), .Q(Q[40]) );
  FD_23 FD_i_41 ( .D(D[41]), .CLK(CLK), .RESET(n16), .Q(Q[41]) );
  FD_22 FD_i_42 ( .D(D[42]), .CLK(CLK), .RESET(n16), .Q(Q[42]) );
  FD_21 FD_i_43 ( .D(D[43]), .CLK(CLK), .RESET(n16), .Q(Q[43]) );
  FD_20 FD_i_44 ( .D(D[44]), .CLK(CLK), .RESET(n16), .Q(Q[44]) );
  FD_19 FD_i_45 ( .D(D[45]), .CLK(CLK), .RESET(n16), .Q(Q[45]) );
  FD_18 FD_i_46 ( .D(D[46]), .CLK(CLK), .RESET(n16), .Q(Q[46]) );
  FD_17 FD_i_47 ( .D(D[47]), .CLK(CLK), .RESET(n17), .Q(Q[47]) );
  FD_16 FD_i_48 ( .D(D[48]), .CLK(CLK), .RESET(n17), .Q(Q[48]) );
  FD_15 FD_i_49 ( .D(D[49]), .CLK(CLK), .RESET(n17), .Q(Q[49]) );
  FD_14 FD_i_50 ( .D(D[50]), .CLK(CLK), .RESET(n16), .Q(Q[50]) );
  FD_13 FD_i_51 ( .D(D[51]), .CLK(CLK), .RESET(n16), .Q(Q[51]) );
  FD_12 FD_i_52 ( .D(D[52]), .CLK(CLK), .RESET(n17), .Q(Q[52]) );
  FD_11 FD_i_53 ( .D(D[53]), .CLK(CLK), .RESET(n16), .Q(Q[53]) );
  FD_10 FD_i_54 ( .D(D[54]), .CLK(CLK), .RESET(n15), .Q(Q[54]) );
  FD_9 FD_i_55 ( .D(D[55]), .CLK(CLK), .RESET(n15), .Q(Q[55]) );
  FD_8 FD_i_56 ( .D(D[56]), .CLK(CLK), .RESET(n15), .Q(Q[56]) );
  FD_7 FD_i_57 ( .D(D[57]), .CLK(CLK), .RESET(n15), .Q(Q[57]) );
  FD_6 FD_i_58 ( .D(D[58]), .CLK(CLK), .RESET(n15), .Q(Q[58]) );
  FD_5 FD_i_59 ( .D(D[59]), .CLK(CLK), .RESET(n15), .Q(Q[59]) );
  FD_4 FD_i_60 ( .D(D[60]), .CLK(CLK), .RESET(n15), .Q(Q[60]) );
  FD_3 FD_i_61 ( .D(D[61]), .CLK(CLK), .RESET(n15), .Q(Q[61]) );
  FD_2 FD_i_62 ( .D(D[62]), .CLK(CLK), .RESET(n15), .Q(Q[62]) );
  FD_1 FD_i_63 ( .D(D[63]), .CLK(CLK), .RESET(n15), .Q(Q[63]) );
  BUF_X1 U1 ( .A(n14), .Z(n19) );
  BUF_X1 U2 ( .A(n14), .Z(n18) );
  BUF_X1 U3 ( .A(n13), .Z(n17) );
  BUF_X1 U4 ( .A(n13), .Z(n16) );
  BUF_X1 U5 ( .A(n13), .Z(n15) );
  BUF_X1 U6 ( .A(n14), .Z(n20) );
  BUF_X1 U7 ( .A(RESET), .Z(n13) );
  BUF_X1 U8 ( .A(RESET), .Z(n14) );
endmodule


module BOOTHMUL_NBIT32 ( INPUT_1, INPUT_2, reset, Clk, MUL_OUT );
  input [31:0] INPUT_1;
  input [31:0] INPUT_2;
  output [63:0] MUL_OUT;
  input reset, Clk;
  wire   \negative_inputs[31][63] , \negative_inputs[31][62] ,
         \negative_inputs[31][61] , \negative_inputs[31][60] ,
         \negative_inputs[31][59] , \negative_inputs[31][58] ,
         \negative_inputs[31][57] , \negative_inputs[31][56] ,
         \negative_inputs[31][55] , \negative_inputs[31][54] ,
         \negative_inputs[31][53] , \negative_inputs[31][52] ,
         \negative_inputs[31][51] , \negative_inputs[31][50] ,
         \negative_inputs[31][49] , \negative_inputs[31][48] ,
         \negative_inputs[31][47] , \negative_inputs[31][46] ,
         \negative_inputs[31][45] , \negative_inputs[31][44] ,
         \negative_inputs[31][43] , \negative_inputs[31][42] ,
         \negative_inputs[31][41] , \negative_inputs[31][40] ,
         \negative_inputs[31][39] , \negative_inputs[31][38] ,
         \negative_inputs[31][37] , \negative_inputs[31][36] ,
         \negative_inputs[31][35] , \negative_inputs[31][34] ,
         \negative_inputs[31][33] , \negative_inputs[31][32] ,
         \negative_inputs[31][31] , \negative_inputs[31][30] ,
         \negative_inputs[31][29] , \negative_inputs[31][28] ,
         \negative_inputs[31][27] , \negative_inputs[31][26] ,
         \negative_inputs[31][25] , \negative_inputs[31][24] ,
         \negative_inputs[31][23] , \negative_inputs[31][22] ,
         \negative_inputs[31][21] , \negative_inputs[31][20] ,
         \negative_inputs[31][19] , \negative_inputs[31][18] ,
         \negative_inputs[31][17] , \negative_inputs[31][16] ,
         \negative_inputs[31][15] , \negative_inputs[31][14] ,
         \negative_inputs[31][13] , \negative_inputs[31][12] ,
         \negative_inputs[31][11] , \negative_inputs[31][10] ,
         \negative_inputs[31][9] , \negative_inputs[31][8] ,
         \negative_inputs[31][7] , \negative_inputs[31][6] ,
         \negative_inputs[31][5] , \negative_inputs[31][4] ,
         \negative_inputs[31][3] , \negative_inputs[31][2] ,
         \negative_inputs[31][1] , \negative_inputs[31][0] ,
         \negative_inputs[30][63] , \negative_inputs[30][62] ,
         \negative_inputs[30][61] , \negative_inputs[30][60] ,
         \negative_inputs[30][59] , \negative_inputs[30][58] ,
         \negative_inputs[30][57] , \negative_inputs[30][56] ,
         \negative_inputs[30][55] , \negative_inputs[30][54] ,
         \negative_inputs[30][53] , \negative_inputs[30][52] ,
         \negative_inputs[30][51] , \negative_inputs[30][50] ,
         \negative_inputs[30][49] , \negative_inputs[30][48] ,
         \negative_inputs[30][47] , \negative_inputs[30][46] ,
         \negative_inputs[30][45] , \negative_inputs[30][44] ,
         \negative_inputs[30][43] , \negative_inputs[30][42] ,
         \negative_inputs[30][41] , \negative_inputs[30][40] ,
         \negative_inputs[30][39] , \negative_inputs[30][38] ,
         \negative_inputs[30][37] , \negative_inputs[30][36] ,
         \negative_inputs[30][35] , \negative_inputs[30][34] ,
         \negative_inputs[30][33] , \negative_inputs[30][32] ,
         \negative_inputs[30][31] , \negative_inputs[30][30] ,
         \negative_inputs[30][29] , \negative_inputs[30][28] ,
         \negative_inputs[30][27] , \negative_inputs[30][26] ,
         \negative_inputs[30][25] , \negative_inputs[30][24] ,
         \negative_inputs[30][23] , \negative_inputs[30][22] ,
         \negative_inputs[30][21] , \negative_inputs[30][20] ,
         \negative_inputs[30][19] , \negative_inputs[30][18] ,
         \negative_inputs[30][17] , \negative_inputs[30][16] ,
         \negative_inputs[30][15] , \negative_inputs[30][14] ,
         \negative_inputs[30][13] , \negative_inputs[30][12] ,
         \negative_inputs[30][11] , \negative_inputs[30][10] ,
         \negative_inputs[30][9] , \negative_inputs[30][8] ,
         \negative_inputs[30][7] , \negative_inputs[30][6] ,
         \negative_inputs[30][5] , \negative_inputs[30][4] ,
         \negative_inputs[30][3] , \negative_inputs[30][2] ,
         \negative_inputs[30][1] , \negative_inputs[30][0] ,
         \negative_inputs[29][63] , \negative_inputs[29][62] ,
         \negative_inputs[29][61] , \negative_inputs[29][60] ,
         \negative_inputs[29][59] , \negative_inputs[29][58] ,
         \negative_inputs[29][57] , \negative_inputs[29][56] ,
         \negative_inputs[29][55] , \negative_inputs[29][54] ,
         \negative_inputs[29][53] , \negative_inputs[29][52] ,
         \negative_inputs[29][51] , \negative_inputs[29][50] ,
         \negative_inputs[29][49] , \negative_inputs[29][48] ,
         \negative_inputs[29][47] , \negative_inputs[29][46] ,
         \negative_inputs[29][45] , \negative_inputs[29][44] ,
         \negative_inputs[29][43] , \negative_inputs[29][42] ,
         \negative_inputs[29][41] , \negative_inputs[29][40] ,
         \negative_inputs[29][39] , \negative_inputs[29][38] ,
         \negative_inputs[29][37] , \negative_inputs[29][36] ,
         \negative_inputs[29][35] , \negative_inputs[29][34] ,
         \negative_inputs[29][33] , \negative_inputs[29][32] ,
         \negative_inputs[29][31] , \negative_inputs[29][30] ,
         \negative_inputs[29][29] , \negative_inputs[29][28] ,
         \negative_inputs[29][27] , \negative_inputs[29][26] ,
         \negative_inputs[29][25] , \negative_inputs[29][24] ,
         \negative_inputs[29][23] , \negative_inputs[29][22] ,
         \negative_inputs[29][21] , \negative_inputs[29][20] ,
         \negative_inputs[29][19] , \negative_inputs[29][18] ,
         \negative_inputs[29][17] , \negative_inputs[29][16] ,
         \negative_inputs[29][15] , \negative_inputs[29][14] ,
         \negative_inputs[29][13] , \negative_inputs[29][12] ,
         \negative_inputs[29][11] , \negative_inputs[29][10] ,
         \negative_inputs[29][9] , \negative_inputs[29][8] ,
         \negative_inputs[29][7] , \negative_inputs[29][6] ,
         \negative_inputs[29][5] , \negative_inputs[29][4] ,
         \negative_inputs[29][3] , \negative_inputs[29][2] ,
         \negative_inputs[29][1] , \negative_inputs[29][0] ,
         \negative_inputs[28][63] , \negative_inputs[28][62] ,
         \negative_inputs[28][61] , \negative_inputs[28][60] ,
         \negative_inputs[28][59] , \negative_inputs[28][58] ,
         \negative_inputs[28][57] , \negative_inputs[28][56] ,
         \negative_inputs[28][55] , \negative_inputs[28][54] ,
         \negative_inputs[28][53] , \negative_inputs[28][52] ,
         \negative_inputs[28][51] , \negative_inputs[28][50] ,
         \negative_inputs[28][49] , \negative_inputs[28][48] ,
         \negative_inputs[28][47] , \negative_inputs[28][46] ,
         \negative_inputs[28][45] , \negative_inputs[28][44] ,
         \negative_inputs[28][43] , \negative_inputs[28][42] ,
         \negative_inputs[28][41] , \negative_inputs[28][40] ,
         \negative_inputs[28][39] , \negative_inputs[28][38] ,
         \negative_inputs[28][37] , \negative_inputs[28][36] ,
         \negative_inputs[28][35] , \negative_inputs[28][34] ,
         \negative_inputs[28][33] , \negative_inputs[28][32] ,
         \negative_inputs[28][31] , \negative_inputs[28][30] ,
         \negative_inputs[28][29] , \negative_inputs[28][28] ,
         \negative_inputs[28][27] , \negative_inputs[28][26] ,
         \negative_inputs[28][25] , \negative_inputs[28][24] ,
         \negative_inputs[28][23] , \negative_inputs[28][22] ,
         \negative_inputs[28][21] , \negative_inputs[28][20] ,
         \negative_inputs[28][19] , \negative_inputs[28][18] ,
         \negative_inputs[28][17] , \negative_inputs[28][16] ,
         \negative_inputs[28][15] , \negative_inputs[28][14] ,
         \negative_inputs[28][13] , \negative_inputs[28][12] ,
         \negative_inputs[28][11] , \negative_inputs[28][10] ,
         \negative_inputs[28][9] , \negative_inputs[28][8] ,
         \negative_inputs[28][7] , \negative_inputs[28][6] ,
         \negative_inputs[28][5] , \negative_inputs[28][4] ,
         \negative_inputs[28][3] , \negative_inputs[28][2] ,
         \negative_inputs[28][1] , \negative_inputs[28][0] ,
         \negative_inputs[27][63] , \negative_inputs[27][62] ,
         \negative_inputs[27][61] , \negative_inputs[27][60] ,
         \negative_inputs[27][59] , \negative_inputs[27][58] ,
         \negative_inputs[27][57] , \negative_inputs[27][56] ,
         \negative_inputs[27][55] , \negative_inputs[27][54] ,
         \negative_inputs[27][53] , \negative_inputs[27][52] ,
         \negative_inputs[27][51] , \negative_inputs[27][50] ,
         \negative_inputs[27][49] , \negative_inputs[27][48] ,
         \negative_inputs[27][47] , \negative_inputs[27][46] ,
         \negative_inputs[27][45] , \negative_inputs[27][44] ,
         \negative_inputs[27][43] , \negative_inputs[27][42] ,
         \negative_inputs[27][41] , \negative_inputs[27][40] ,
         \negative_inputs[27][39] , \negative_inputs[27][38] ,
         \negative_inputs[27][37] , \negative_inputs[27][36] ,
         \negative_inputs[27][35] , \negative_inputs[27][34] ,
         \negative_inputs[27][33] , \negative_inputs[27][32] ,
         \negative_inputs[27][31] , \negative_inputs[27][30] ,
         \negative_inputs[27][29] , \negative_inputs[27][28] ,
         \negative_inputs[27][27] , \negative_inputs[27][26] ,
         \negative_inputs[27][25] , \negative_inputs[27][24] ,
         \negative_inputs[27][23] , \negative_inputs[27][22] ,
         \negative_inputs[27][21] , \negative_inputs[27][20] ,
         \negative_inputs[27][19] , \negative_inputs[27][18] ,
         \negative_inputs[27][17] , \negative_inputs[27][16] ,
         \negative_inputs[27][15] , \negative_inputs[27][14] ,
         \negative_inputs[27][13] , \negative_inputs[27][12] ,
         \negative_inputs[27][11] , \negative_inputs[27][10] ,
         \negative_inputs[27][9] , \negative_inputs[27][8] ,
         \negative_inputs[27][7] , \negative_inputs[27][6] ,
         \negative_inputs[27][5] , \negative_inputs[27][4] ,
         \negative_inputs[27][3] , \negative_inputs[27][2] ,
         \negative_inputs[27][1] , \negative_inputs[27][0] ,
         \negative_inputs[26][63] , \negative_inputs[26][62] ,
         \negative_inputs[26][61] , \negative_inputs[26][60] ,
         \negative_inputs[26][59] , \negative_inputs[26][58] ,
         \negative_inputs[26][57] , \negative_inputs[26][56] ,
         \negative_inputs[26][55] , \negative_inputs[26][54] ,
         \negative_inputs[26][53] , \negative_inputs[26][52] ,
         \negative_inputs[26][51] , \negative_inputs[26][50] ,
         \negative_inputs[26][49] , \negative_inputs[26][48] ,
         \negative_inputs[26][47] , \negative_inputs[26][46] ,
         \negative_inputs[26][45] , \negative_inputs[26][44] ,
         \negative_inputs[26][43] , \negative_inputs[26][42] ,
         \negative_inputs[26][41] , \negative_inputs[26][40] ,
         \negative_inputs[26][39] , \negative_inputs[26][38] ,
         \negative_inputs[26][37] , \negative_inputs[26][36] ,
         \negative_inputs[26][35] , \negative_inputs[26][34] ,
         \negative_inputs[26][33] , \negative_inputs[26][32] ,
         \negative_inputs[26][31] , \negative_inputs[26][30] ,
         \negative_inputs[26][29] , \negative_inputs[26][28] ,
         \negative_inputs[26][27] , \negative_inputs[26][26] ,
         \negative_inputs[26][25] , \negative_inputs[26][24] ,
         \negative_inputs[26][23] , \negative_inputs[26][22] ,
         \negative_inputs[26][21] , \negative_inputs[26][20] ,
         \negative_inputs[26][19] , \negative_inputs[26][18] ,
         \negative_inputs[26][17] , \negative_inputs[26][16] ,
         \negative_inputs[26][15] , \negative_inputs[26][14] ,
         \negative_inputs[26][13] , \negative_inputs[26][12] ,
         \negative_inputs[26][11] , \negative_inputs[26][10] ,
         \negative_inputs[26][9] , \negative_inputs[26][8] ,
         \negative_inputs[26][7] , \negative_inputs[26][6] ,
         \negative_inputs[26][5] , \negative_inputs[26][4] ,
         \negative_inputs[26][3] , \negative_inputs[26][2] ,
         \negative_inputs[26][1] , \negative_inputs[26][0] ,
         \negative_inputs[25][63] , \negative_inputs[25][62] ,
         \negative_inputs[25][61] , \negative_inputs[25][60] ,
         \negative_inputs[25][59] , \negative_inputs[25][58] ,
         \negative_inputs[25][57] , \negative_inputs[25][56] ,
         \negative_inputs[25][55] , \negative_inputs[25][54] ,
         \negative_inputs[25][53] , \negative_inputs[25][52] ,
         \negative_inputs[25][51] , \negative_inputs[25][50] ,
         \negative_inputs[25][49] , \negative_inputs[25][48] ,
         \negative_inputs[25][47] , \negative_inputs[25][46] ,
         \negative_inputs[25][45] , \negative_inputs[25][44] ,
         \negative_inputs[25][43] , \negative_inputs[25][42] ,
         \negative_inputs[25][41] , \negative_inputs[25][40] ,
         \negative_inputs[25][39] , \negative_inputs[25][38] ,
         \negative_inputs[25][37] , \negative_inputs[25][36] ,
         \negative_inputs[25][35] , \negative_inputs[25][34] ,
         \negative_inputs[25][33] , \negative_inputs[25][32] ,
         \negative_inputs[25][31] , \negative_inputs[25][30] ,
         \negative_inputs[25][29] , \negative_inputs[25][28] ,
         \negative_inputs[25][27] , \negative_inputs[25][26] ,
         \negative_inputs[25][25] , \negative_inputs[25][24] ,
         \negative_inputs[25][23] , \negative_inputs[25][22] ,
         \negative_inputs[25][21] , \negative_inputs[25][20] ,
         \negative_inputs[25][19] , \negative_inputs[25][18] ,
         \negative_inputs[25][17] , \negative_inputs[25][16] ,
         \negative_inputs[25][15] , \negative_inputs[25][14] ,
         \negative_inputs[25][13] , \negative_inputs[25][12] ,
         \negative_inputs[25][11] , \negative_inputs[25][10] ,
         \negative_inputs[25][9] , \negative_inputs[25][8] ,
         \negative_inputs[25][7] , \negative_inputs[25][6] ,
         \negative_inputs[25][5] , \negative_inputs[25][4] ,
         \negative_inputs[25][3] , \negative_inputs[25][2] ,
         \negative_inputs[25][1] , \negative_inputs[25][0] ,
         \negative_inputs[24][63] , \negative_inputs[24][62] ,
         \negative_inputs[24][61] , \negative_inputs[24][60] ,
         \negative_inputs[24][59] , \negative_inputs[24][58] ,
         \negative_inputs[24][57] , \negative_inputs[24][56] ,
         \negative_inputs[24][55] , \negative_inputs[24][54] ,
         \negative_inputs[24][53] , \negative_inputs[24][52] ,
         \negative_inputs[24][51] , \negative_inputs[24][50] ,
         \negative_inputs[24][49] , \negative_inputs[24][48] ,
         \negative_inputs[24][47] , \negative_inputs[24][46] ,
         \negative_inputs[24][45] , \negative_inputs[24][44] ,
         \negative_inputs[24][43] , \negative_inputs[24][42] ,
         \negative_inputs[24][41] , \negative_inputs[24][40] ,
         \negative_inputs[24][39] , \negative_inputs[24][38] ,
         \negative_inputs[24][37] , \negative_inputs[24][36] ,
         \negative_inputs[24][35] , \negative_inputs[24][34] ,
         \negative_inputs[24][33] , \negative_inputs[24][32] ,
         \negative_inputs[24][31] , \negative_inputs[24][30] ,
         \negative_inputs[24][29] , \negative_inputs[24][28] ,
         \negative_inputs[24][27] , \negative_inputs[24][26] ,
         \negative_inputs[24][25] , \negative_inputs[24][24] ,
         \negative_inputs[24][23] , \negative_inputs[24][22] ,
         \negative_inputs[24][21] , \negative_inputs[24][20] ,
         \negative_inputs[24][19] , \negative_inputs[24][18] ,
         \negative_inputs[24][17] , \negative_inputs[24][16] ,
         \negative_inputs[24][15] , \negative_inputs[24][14] ,
         \negative_inputs[24][13] , \negative_inputs[24][12] ,
         \negative_inputs[24][11] , \negative_inputs[24][10] ,
         \negative_inputs[24][9] , \negative_inputs[24][8] ,
         \negative_inputs[24][7] , \negative_inputs[24][6] ,
         \negative_inputs[24][5] , \negative_inputs[24][4] ,
         \negative_inputs[24][3] , \negative_inputs[24][2] ,
         \negative_inputs[24][1] , \negative_inputs[24][0] ,
         \negative_inputs[23][63] , \negative_inputs[23][62] ,
         \negative_inputs[23][61] , \negative_inputs[23][60] ,
         \negative_inputs[23][59] , \negative_inputs[23][58] ,
         \negative_inputs[23][57] , \negative_inputs[23][56] ,
         \negative_inputs[23][55] , \negative_inputs[23][54] ,
         \negative_inputs[23][53] , \negative_inputs[23][52] ,
         \negative_inputs[23][51] , \negative_inputs[23][50] ,
         \negative_inputs[23][49] , \negative_inputs[23][48] ,
         \negative_inputs[23][47] , \negative_inputs[23][46] ,
         \negative_inputs[23][45] , \negative_inputs[23][44] ,
         \negative_inputs[23][43] , \negative_inputs[23][42] ,
         \negative_inputs[23][41] , \negative_inputs[23][40] ,
         \negative_inputs[23][39] , \negative_inputs[23][38] ,
         \negative_inputs[23][37] , \negative_inputs[23][36] ,
         \negative_inputs[23][35] , \negative_inputs[23][34] ,
         \negative_inputs[23][33] , \negative_inputs[23][32] ,
         \negative_inputs[23][31] , \negative_inputs[23][30] ,
         \negative_inputs[23][29] , \negative_inputs[23][28] ,
         \negative_inputs[23][27] , \negative_inputs[23][26] ,
         \negative_inputs[23][25] , \negative_inputs[23][24] ,
         \negative_inputs[23][23] , \negative_inputs[23][22] ,
         \negative_inputs[23][21] , \negative_inputs[23][20] ,
         \negative_inputs[23][19] , \negative_inputs[23][18] ,
         \negative_inputs[23][17] , \negative_inputs[23][16] ,
         \negative_inputs[23][15] , \negative_inputs[23][14] ,
         \negative_inputs[23][13] , \negative_inputs[23][12] ,
         \negative_inputs[23][11] , \negative_inputs[23][10] ,
         \negative_inputs[23][9] , \negative_inputs[23][8] ,
         \negative_inputs[23][7] , \negative_inputs[23][6] ,
         \negative_inputs[23][5] , \negative_inputs[23][4] ,
         \negative_inputs[23][3] , \negative_inputs[23][2] ,
         \negative_inputs[23][1] , \negative_inputs[23][0] ,
         \negative_inputs[22][63] , \negative_inputs[22][62] ,
         \negative_inputs[22][61] , \negative_inputs[22][60] ,
         \negative_inputs[22][59] , \negative_inputs[22][58] ,
         \negative_inputs[22][57] , \negative_inputs[22][56] ,
         \negative_inputs[22][55] , \negative_inputs[22][54] ,
         \negative_inputs[22][53] , \negative_inputs[22][52] ,
         \negative_inputs[22][51] , \negative_inputs[22][50] ,
         \negative_inputs[22][49] , \negative_inputs[22][48] ,
         \negative_inputs[22][47] , \negative_inputs[22][46] ,
         \negative_inputs[22][45] , \negative_inputs[22][44] ,
         \negative_inputs[22][43] , \negative_inputs[22][42] ,
         \negative_inputs[22][41] , \negative_inputs[22][40] ,
         \negative_inputs[22][39] , \negative_inputs[22][38] ,
         \negative_inputs[22][37] , \negative_inputs[22][36] ,
         \negative_inputs[22][35] , \negative_inputs[22][34] ,
         \negative_inputs[22][33] , \negative_inputs[22][32] ,
         \negative_inputs[22][31] , \negative_inputs[22][30] ,
         \negative_inputs[22][29] , \negative_inputs[22][28] ,
         \negative_inputs[22][27] , \negative_inputs[22][26] ,
         \negative_inputs[22][25] , \negative_inputs[22][24] ,
         \negative_inputs[22][23] , \negative_inputs[22][22] ,
         \negative_inputs[22][21] , \negative_inputs[22][20] ,
         \negative_inputs[22][19] , \negative_inputs[22][18] ,
         \negative_inputs[22][17] , \negative_inputs[22][16] ,
         \negative_inputs[22][15] , \negative_inputs[22][14] ,
         \negative_inputs[22][13] , \negative_inputs[22][12] ,
         \negative_inputs[22][11] , \negative_inputs[22][10] ,
         \negative_inputs[22][9] , \negative_inputs[22][8] ,
         \negative_inputs[22][7] , \negative_inputs[22][6] ,
         \negative_inputs[22][5] , \negative_inputs[22][4] ,
         \negative_inputs[22][3] , \negative_inputs[22][2] ,
         \negative_inputs[22][1] , \negative_inputs[22][0] ,
         \negative_inputs[21][63] , \negative_inputs[21][62] ,
         \negative_inputs[21][61] , \negative_inputs[21][60] ,
         \negative_inputs[21][59] , \negative_inputs[21][58] ,
         \negative_inputs[21][57] , \negative_inputs[21][56] ,
         \negative_inputs[21][55] , \negative_inputs[21][54] ,
         \negative_inputs[21][53] , \negative_inputs[21][52] ,
         \negative_inputs[21][51] , \negative_inputs[21][50] ,
         \negative_inputs[21][49] , \negative_inputs[21][48] ,
         \negative_inputs[21][47] , \negative_inputs[21][46] ,
         \negative_inputs[21][45] , \negative_inputs[21][44] ,
         \negative_inputs[21][43] , \negative_inputs[21][42] ,
         \negative_inputs[21][41] , \negative_inputs[21][40] ,
         \negative_inputs[21][39] , \negative_inputs[21][38] ,
         \negative_inputs[21][37] , \negative_inputs[21][36] ,
         \negative_inputs[21][35] , \negative_inputs[21][34] ,
         \negative_inputs[21][33] , \negative_inputs[21][32] ,
         \negative_inputs[21][31] , \negative_inputs[21][30] ,
         \negative_inputs[21][29] , \negative_inputs[21][28] ,
         \negative_inputs[21][27] , \negative_inputs[21][26] ,
         \negative_inputs[21][25] , \negative_inputs[21][24] ,
         \negative_inputs[21][23] , \negative_inputs[21][22] ,
         \negative_inputs[21][21] , \negative_inputs[21][20] ,
         \negative_inputs[21][19] , \negative_inputs[21][18] ,
         \negative_inputs[21][17] , \negative_inputs[21][16] ,
         \negative_inputs[21][15] , \negative_inputs[21][14] ,
         \negative_inputs[21][13] , \negative_inputs[21][12] ,
         \negative_inputs[21][11] , \negative_inputs[21][10] ,
         \negative_inputs[21][9] , \negative_inputs[21][8] ,
         \negative_inputs[21][7] , \negative_inputs[21][6] ,
         \negative_inputs[21][5] , \negative_inputs[21][4] ,
         \negative_inputs[21][3] , \negative_inputs[21][2] ,
         \negative_inputs[21][1] , \negative_inputs[21][0] ,
         \negative_inputs[20][63] , \negative_inputs[20][62] ,
         \negative_inputs[20][61] , \negative_inputs[20][60] ,
         \negative_inputs[20][59] , \negative_inputs[20][58] ,
         \negative_inputs[20][57] , \negative_inputs[20][56] ,
         \negative_inputs[20][55] , \negative_inputs[20][54] ,
         \negative_inputs[20][53] , \negative_inputs[20][52] ,
         \negative_inputs[20][51] , \negative_inputs[20][50] ,
         \negative_inputs[20][49] , \negative_inputs[20][48] ,
         \negative_inputs[20][47] , \negative_inputs[20][46] ,
         \negative_inputs[20][45] , \negative_inputs[20][44] ,
         \negative_inputs[20][43] , \negative_inputs[20][42] ,
         \negative_inputs[20][41] , \negative_inputs[20][40] ,
         \negative_inputs[20][39] , \negative_inputs[20][38] ,
         \negative_inputs[20][37] , \negative_inputs[20][36] ,
         \negative_inputs[20][35] , \negative_inputs[20][34] ,
         \negative_inputs[20][33] , \negative_inputs[20][32] ,
         \negative_inputs[20][31] , \negative_inputs[20][30] ,
         \negative_inputs[20][29] , \negative_inputs[20][28] ,
         \negative_inputs[20][27] , \negative_inputs[20][26] ,
         \negative_inputs[20][25] , \negative_inputs[20][24] ,
         \negative_inputs[20][23] , \negative_inputs[20][22] ,
         \negative_inputs[20][21] , \negative_inputs[20][20] ,
         \negative_inputs[20][19] , \negative_inputs[20][18] ,
         \negative_inputs[20][17] , \negative_inputs[20][16] ,
         \negative_inputs[20][15] , \negative_inputs[20][14] ,
         \negative_inputs[20][13] , \negative_inputs[20][12] ,
         \negative_inputs[20][11] , \negative_inputs[20][10] ,
         \negative_inputs[20][9] , \negative_inputs[20][8] ,
         \negative_inputs[20][7] , \negative_inputs[20][6] ,
         \negative_inputs[20][5] , \negative_inputs[20][4] ,
         \negative_inputs[20][3] , \negative_inputs[20][2] ,
         \negative_inputs[20][1] , \negative_inputs[20][0] ,
         \negative_inputs[19][63] , \negative_inputs[19][62] ,
         \negative_inputs[19][61] , \negative_inputs[19][60] ,
         \negative_inputs[19][59] , \negative_inputs[19][58] ,
         \negative_inputs[19][57] , \negative_inputs[19][56] ,
         \negative_inputs[19][55] , \negative_inputs[19][54] ,
         \negative_inputs[19][53] , \negative_inputs[19][52] ,
         \negative_inputs[19][51] , \negative_inputs[19][50] ,
         \negative_inputs[19][49] , \negative_inputs[19][48] ,
         \negative_inputs[19][47] , \negative_inputs[19][46] ,
         \negative_inputs[19][45] , \negative_inputs[19][44] ,
         \negative_inputs[19][43] , \negative_inputs[19][42] ,
         \negative_inputs[19][41] , \negative_inputs[19][40] ,
         \negative_inputs[19][39] , \negative_inputs[19][38] ,
         \negative_inputs[19][37] , \negative_inputs[19][36] ,
         \negative_inputs[19][35] , \negative_inputs[19][34] ,
         \negative_inputs[19][33] , \negative_inputs[19][32] ,
         \negative_inputs[19][31] , \negative_inputs[19][30] ,
         \negative_inputs[19][29] , \negative_inputs[19][28] ,
         \negative_inputs[19][27] , \negative_inputs[19][26] ,
         \negative_inputs[19][25] , \negative_inputs[19][24] ,
         \negative_inputs[19][23] , \negative_inputs[19][22] ,
         \negative_inputs[19][21] , \negative_inputs[19][20] ,
         \negative_inputs[19][19] , \negative_inputs[19][18] ,
         \negative_inputs[19][17] , \negative_inputs[19][16] ,
         \negative_inputs[19][15] , \negative_inputs[19][14] ,
         \negative_inputs[19][13] , \negative_inputs[19][12] ,
         \negative_inputs[19][11] , \negative_inputs[19][10] ,
         \negative_inputs[19][9] , \negative_inputs[19][8] ,
         \negative_inputs[19][7] , \negative_inputs[19][6] ,
         \negative_inputs[19][5] , \negative_inputs[19][4] ,
         \negative_inputs[19][3] , \negative_inputs[19][2] ,
         \negative_inputs[19][1] , \negative_inputs[19][0] ,
         \negative_inputs[18][63] , \negative_inputs[18][62] ,
         \negative_inputs[18][61] , \negative_inputs[18][60] ,
         \negative_inputs[18][59] , \negative_inputs[18][58] ,
         \negative_inputs[18][57] , \negative_inputs[18][56] ,
         \negative_inputs[18][55] , \negative_inputs[18][54] ,
         \negative_inputs[18][53] , \negative_inputs[18][52] ,
         \negative_inputs[18][51] , \negative_inputs[18][50] ,
         \negative_inputs[18][49] , \negative_inputs[18][48] ,
         \negative_inputs[18][47] , \negative_inputs[18][46] ,
         \negative_inputs[18][45] , \negative_inputs[18][44] ,
         \negative_inputs[18][43] , \negative_inputs[18][42] ,
         \negative_inputs[18][41] , \negative_inputs[18][40] ,
         \negative_inputs[18][39] , \negative_inputs[18][38] ,
         \negative_inputs[18][37] , \negative_inputs[18][36] ,
         \negative_inputs[18][35] , \negative_inputs[18][34] ,
         \negative_inputs[18][33] , \negative_inputs[18][32] ,
         \negative_inputs[18][31] , \negative_inputs[18][30] ,
         \negative_inputs[18][29] , \negative_inputs[18][28] ,
         \negative_inputs[18][27] , \negative_inputs[18][26] ,
         \negative_inputs[18][25] , \negative_inputs[18][24] ,
         \negative_inputs[18][23] , \negative_inputs[18][22] ,
         \negative_inputs[18][21] , \negative_inputs[18][20] ,
         \negative_inputs[18][19] , \negative_inputs[18][18] ,
         \negative_inputs[18][17] , \negative_inputs[18][16] ,
         \negative_inputs[18][15] , \negative_inputs[18][14] ,
         \negative_inputs[18][13] , \negative_inputs[18][12] ,
         \negative_inputs[18][11] , \negative_inputs[18][10] ,
         \negative_inputs[18][9] , \negative_inputs[18][8] ,
         \negative_inputs[18][7] , \negative_inputs[18][6] ,
         \negative_inputs[18][5] , \negative_inputs[18][4] ,
         \negative_inputs[18][3] , \negative_inputs[18][2] ,
         \negative_inputs[18][1] , \negative_inputs[18][0] ,
         \negative_inputs[17][63] , \negative_inputs[17][62] ,
         \negative_inputs[17][61] , \negative_inputs[17][60] ,
         \negative_inputs[17][59] , \negative_inputs[17][58] ,
         \negative_inputs[17][57] , \negative_inputs[17][56] ,
         \negative_inputs[17][55] , \negative_inputs[17][54] ,
         \negative_inputs[17][53] , \negative_inputs[17][52] ,
         \negative_inputs[17][51] , \negative_inputs[17][50] ,
         \negative_inputs[17][49] , \negative_inputs[17][48] ,
         \negative_inputs[17][47] , \negative_inputs[17][46] ,
         \negative_inputs[17][45] , \negative_inputs[17][44] ,
         \negative_inputs[17][43] , \negative_inputs[17][42] ,
         \negative_inputs[17][41] , \negative_inputs[17][40] ,
         \negative_inputs[17][39] , \negative_inputs[17][38] ,
         \negative_inputs[17][37] , \negative_inputs[17][36] ,
         \negative_inputs[17][35] , \negative_inputs[17][34] ,
         \negative_inputs[17][33] , \negative_inputs[17][32] ,
         \negative_inputs[17][31] , \negative_inputs[17][30] ,
         \negative_inputs[17][29] , \negative_inputs[17][28] ,
         \negative_inputs[17][27] , \negative_inputs[17][26] ,
         \negative_inputs[17][25] , \negative_inputs[17][24] ,
         \negative_inputs[17][23] , \negative_inputs[17][22] ,
         \negative_inputs[17][21] , \negative_inputs[17][20] ,
         \negative_inputs[17][19] , \negative_inputs[17][18] ,
         \negative_inputs[17][17] , \negative_inputs[17][16] ,
         \negative_inputs[17][15] , \negative_inputs[17][14] ,
         \negative_inputs[17][13] , \negative_inputs[17][12] ,
         \negative_inputs[17][11] , \negative_inputs[17][10] ,
         \negative_inputs[17][9] , \negative_inputs[17][8] ,
         \negative_inputs[17][7] , \negative_inputs[17][6] ,
         \negative_inputs[17][5] , \negative_inputs[17][4] ,
         \negative_inputs[17][3] , \negative_inputs[17][2] ,
         \negative_inputs[17][1] , \negative_inputs[17][0] ,
         \negative_inputs[16][63] , \negative_inputs[16][62] ,
         \negative_inputs[16][61] , \negative_inputs[16][60] ,
         \negative_inputs[16][59] , \negative_inputs[16][58] ,
         \negative_inputs[16][57] , \negative_inputs[16][56] ,
         \negative_inputs[16][55] , \negative_inputs[16][54] ,
         \negative_inputs[16][53] , \negative_inputs[16][52] ,
         \negative_inputs[16][51] , \negative_inputs[16][50] ,
         \negative_inputs[16][49] , \negative_inputs[16][48] ,
         \negative_inputs[16][47] , \negative_inputs[16][46] ,
         \negative_inputs[16][45] , \negative_inputs[16][44] ,
         \negative_inputs[16][43] , \negative_inputs[16][42] ,
         \negative_inputs[16][41] , \negative_inputs[16][40] ,
         \negative_inputs[16][39] , \negative_inputs[16][38] ,
         \negative_inputs[16][37] , \negative_inputs[16][36] ,
         \negative_inputs[16][35] , \negative_inputs[16][34] ,
         \negative_inputs[16][33] , \negative_inputs[16][32] ,
         \negative_inputs[16][31] , \negative_inputs[16][30] ,
         \negative_inputs[16][29] , \negative_inputs[16][28] ,
         \negative_inputs[16][27] , \negative_inputs[16][26] ,
         \negative_inputs[16][25] , \negative_inputs[16][24] ,
         \negative_inputs[16][23] , \negative_inputs[16][22] ,
         \negative_inputs[16][21] , \negative_inputs[16][20] ,
         \negative_inputs[16][19] , \negative_inputs[16][18] ,
         \negative_inputs[16][17] , \negative_inputs[16][16] ,
         \negative_inputs[16][15] , \negative_inputs[16][14] ,
         \negative_inputs[16][13] , \negative_inputs[16][12] ,
         \negative_inputs[16][11] , \negative_inputs[16][10] ,
         \negative_inputs[16][9] , \negative_inputs[16][8] ,
         \negative_inputs[16][7] , \negative_inputs[16][6] ,
         \negative_inputs[16][5] , \negative_inputs[16][4] ,
         \negative_inputs[16][3] , \negative_inputs[16][2] ,
         \negative_inputs[16][1] , \negative_inputs[16][0] ,
         \negative_inputs[15][63] , \negative_inputs[15][62] ,
         \negative_inputs[15][61] , \negative_inputs[15][60] ,
         \negative_inputs[15][59] , \negative_inputs[15][58] ,
         \negative_inputs[15][57] , \negative_inputs[15][56] ,
         \negative_inputs[15][55] , \negative_inputs[15][54] ,
         \negative_inputs[15][53] , \negative_inputs[15][52] ,
         \negative_inputs[15][51] , \negative_inputs[15][50] ,
         \negative_inputs[15][49] , \negative_inputs[15][48] ,
         \negative_inputs[15][47] , \negative_inputs[15][46] ,
         \negative_inputs[15][45] , \negative_inputs[15][44] ,
         \negative_inputs[15][43] , \negative_inputs[15][42] ,
         \negative_inputs[15][41] , \negative_inputs[15][40] ,
         \negative_inputs[15][39] , \negative_inputs[15][38] ,
         \negative_inputs[15][37] , \negative_inputs[15][36] ,
         \negative_inputs[15][35] , \negative_inputs[15][34] ,
         \negative_inputs[15][33] , \negative_inputs[15][32] ,
         \negative_inputs[15][31] , \negative_inputs[15][30] ,
         \negative_inputs[15][29] , \negative_inputs[15][28] ,
         \negative_inputs[15][27] , \negative_inputs[15][26] ,
         \negative_inputs[15][25] , \negative_inputs[15][24] ,
         \negative_inputs[15][23] , \negative_inputs[15][22] ,
         \negative_inputs[15][21] , \negative_inputs[15][20] ,
         \negative_inputs[15][19] , \negative_inputs[15][18] ,
         \negative_inputs[15][17] , \negative_inputs[15][16] ,
         \negative_inputs[15][15] , \negative_inputs[15][14] ,
         \negative_inputs[15][13] , \negative_inputs[15][12] ,
         \negative_inputs[15][11] , \negative_inputs[15][10] ,
         \negative_inputs[15][9] , \negative_inputs[15][8] ,
         \negative_inputs[15][7] , \negative_inputs[15][6] ,
         \negative_inputs[15][5] , \negative_inputs[15][4] ,
         \negative_inputs[15][3] , \negative_inputs[15][2] ,
         \negative_inputs[15][1] , \negative_inputs[15][0] ,
         \negative_inputs[14][63] , \negative_inputs[14][62] ,
         \negative_inputs[14][61] , \negative_inputs[14][60] ,
         \negative_inputs[14][59] , \negative_inputs[14][58] ,
         \negative_inputs[14][57] , \negative_inputs[14][56] ,
         \negative_inputs[14][55] , \negative_inputs[14][54] ,
         \negative_inputs[14][53] , \negative_inputs[14][52] ,
         \negative_inputs[14][51] , \negative_inputs[14][50] ,
         \negative_inputs[14][49] , \negative_inputs[14][48] ,
         \negative_inputs[14][47] , \negative_inputs[14][46] ,
         \negative_inputs[14][45] , \negative_inputs[14][44] ,
         \negative_inputs[14][43] , \negative_inputs[14][42] ,
         \negative_inputs[14][41] , \negative_inputs[14][40] ,
         \negative_inputs[14][39] , \negative_inputs[14][38] ,
         \negative_inputs[14][37] , \negative_inputs[14][36] ,
         \negative_inputs[14][35] , \negative_inputs[14][34] ,
         \negative_inputs[14][33] , \negative_inputs[14][32] ,
         \negative_inputs[14][31] , \negative_inputs[14][30] ,
         \negative_inputs[14][29] , \negative_inputs[14][28] ,
         \negative_inputs[14][27] , \negative_inputs[14][26] ,
         \negative_inputs[14][25] , \negative_inputs[14][24] ,
         \negative_inputs[14][23] , \negative_inputs[14][22] ,
         \negative_inputs[14][21] , \negative_inputs[14][20] ,
         \negative_inputs[14][19] , \negative_inputs[14][18] ,
         \negative_inputs[14][17] , \negative_inputs[14][16] ,
         \negative_inputs[14][15] , \negative_inputs[14][14] ,
         \negative_inputs[14][13] , \negative_inputs[14][12] ,
         \negative_inputs[14][11] , \negative_inputs[14][10] ,
         \negative_inputs[14][9] , \negative_inputs[14][8] ,
         \negative_inputs[14][7] , \negative_inputs[14][6] ,
         \negative_inputs[14][5] , \negative_inputs[14][4] ,
         \negative_inputs[14][3] , \negative_inputs[14][2] ,
         \negative_inputs[14][1] , \negative_inputs[14][0] ,
         \negative_inputs[13][63] , \negative_inputs[13][62] ,
         \negative_inputs[13][61] , \negative_inputs[13][60] ,
         \negative_inputs[13][59] , \negative_inputs[13][58] ,
         \negative_inputs[13][57] , \negative_inputs[13][56] ,
         \negative_inputs[13][55] , \negative_inputs[13][54] ,
         \negative_inputs[13][53] , \negative_inputs[13][52] ,
         \negative_inputs[13][51] , \negative_inputs[13][50] ,
         \negative_inputs[13][49] , \negative_inputs[13][48] ,
         \negative_inputs[13][47] , \negative_inputs[13][46] ,
         \negative_inputs[13][45] , \negative_inputs[13][44] ,
         \negative_inputs[13][43] , \negative_inputs[13][42] ,
         \negative_inputs[13][41] , \negative_inputs[13][40] ,
         \negative_inputs[13][39] , \negative_inputs[13][38] ,
         \negative_inputs[13][37] , \negative_inputs[13][36] ,
         \negative_inputs[13][35] , \negative_inputs[13][34] ,
         \negative_inputs[13][33] , \negative_inputs[13][32] ,
         \negative_inputs[13][31] , \negative_inputs[13][30] ,
         \negative_inputs[13][29] , \negative_inputs[13][28] ,
         \negative_inputs[13][27] , \negative_inputs[13][26] ,
         \negative_inputs[13][25] , \negative_inputs[13][24] ,
         \negative_inputs[13][23] , \negative_inputs[13][22] ,
         \negative_inputs[13][21] , \negative_inputs[13][20] ,
         \negative_inputs[13][19] , \negative_inputs[13][18] ,
         \negative_inputs[13][17] , \negative_inputs[13][16] ,
         \negative_inputs[13][15] , \negative_inputs[13][14] ,
         \negative_inputs[13][13] , \negative_inputs[13][12] ,
         \negative_inputs[13][11] , \negative_inputs[13][10] ,
         \negative_inputs[13][9] , \negative_inputs[13][8] ,
         \negative_inputs[13][7] , \negative_inputs[13][6] ,
         \negative_inputs[13][5] , \negative_inputs[13][4] ,
         \negative_inputs[13][3] , \negative_inputs[13][2] ,
         \negative_inputs[13][1] , \negative_inputs[13][0] ,
         \negative_inputs[12][63] , \negative_inputs[12][62] ,
         \negative_inputs[12][61] , \negative_inputs[12][60] ,
         \negative_inputs[12][59] , \negative_inputs[12][58] ,
         \negative_inputs[12][57] , \negative_inputs[12][56] ,
         \negative_inputs[12][55] , \negative_inputs[12][54] ,
         \negative_inputs[12][53] , \negative_inputs[12][52] ,
         \negative_inputs[12][51] , \negative_inputs[12][50] ,
         \negative_inputs[12][49] , \negative_inputs[12][48] ,
         \negative_inputs[12][47] , \negative_inputs[12][46] ,
         \negative_inputs[12][45] , \negative_inputs[12][44] ,
         \negative_inputs[12][43] , \negative_inputs[12][42] ,
         \negative_inputs[12][41] , \negative_inputs[12][40] ,
         \negative_inputs[12][39] , \negative_inputs[12][38] ,
         \negative_inputs[12][37] , \negative_inputs[12][36] ,
         \negative_inputs[12][35] , \negative_inputs[12][34] ,
         \negative_inputs[12][33] , \negative_inputs[12][32] ,
         \negative_inputs[12][31] , \negative_inputs[12][30] ,
         \negative_inputs[12][29] , \negative_inputs[12][28] ,
         \negative_inputs[12][27] , \negative_inputs[12][26] ,
         \negative_inputs[12][25] , \negative_inputs[12][24] ,
         \negative_inputs[12][23] , \negative_inputs[12][22] ,
         \negative_inputs[12][21] , \negative_inputs[12][20] ,
         \negative_inputs[12][19] , \negative_inputs[12][18] ,
         \negative_inputs[12][17] , \negative_inputs[12][16] ,
         \negative_inputs[12][15] , \negative_inputs[12][14] ,
         \negative_inputs[12][13] , \negative_inputs[12][12] ,
         \negative_inputs[12][11] , \negative_inputs[12][10] ,
         \negative_inputs[12][9] , \negative_inputs[12][8] ,
         \negative_inputs[12][7] , \negative_inputs[12][6] ,
         \negative_inputs[12][5] , \negative_inputs[12][4] ,
         \negative_inputs[12][3] , \negative_inputs[12][2] ,
         \negative_inputs[12][1] , \negative_inputs[12][0] ,
         \negative_inputs[11][63] , \negative_inputs[11][62] ,
         \negative_inputs[11][61] , \negative_inputs[11][60] ,
         \negative_inputs[11][59] , \negative_inputs[11][58] ,
         \negative_inputs[11][57] , \negative_inputs[11][56] ,
         \negative_inputs[11][55] , \negative_inputs[11][54] ,
         \negative_inputs[11][53] , \negative_inputs[11][52] ,
         \negative_inputs[11][51] , \negative_inputs[11][50] ,
         \negative_inputs[11][49] , \negative_inputs[11][48] ,
         \negative_inputs[11][47] , \negative_inputs[11][46] ,
         \negative_inputs[11][45] , \negative_inputs[11][44] ,
         \negative_inputs[11][43] , \negative_inputs[11][42] ,
         \negative_inputs[11][41] , \negative_inputs[11][40] ,
         \negative_inputs[11][39] , \negative_inputs[11][38] ,
         \negative_inputs[11][37] , \negative_inputs[11][36] ,
         \negative_inputs[11][35] , \negative_inputs[11][34] ,
         \negative_inputs[11][33] , \negative_inputs[11][32] ,
         \negative_inputs[11][31] , \negative_inputs[11][30] ,
         \negative_inputs[11][29] , \negative_inputs[11][28] ,
         \negative_inputs[11][27] , \negative_inputs[11][26] ,
         \negative_inputs[11][25] , \negative_inputs[11][24] ,
         \negative_inputs[11][23] , \negative_inputs[11][22] ,
         \negative_inputs[11][21] , \negative_inputs[11][20] ,
         \negative_inputs[11][19] , \negative_inputs[11][18] ,
         \negative_inputs[11][17] , \negative_inputs[11][16] ,
         \negative_inputs[11][15] , \negative_inputs[11][14] ,
         \negative_inputs[11][13] , \negative_inputs[11][12] ,
         \negative_inputs[11][11] , \negative_inputs[11][10] ,
         \negative_inputs[11][9] , \negative_inputs[11][8] ,
         \negative_inputs[11][7] , \negative_inputs[11][6] ,
         \negative_inputs[11][5] , \negative_inputs[11][4] ,
         \negative_inputs[11][3] , \negative_inputs[11][2] ,
         \negative_inputs[11][1] , \negative_inputs[11][0] ,
         \negative_inputs[10][63] , \negative_inputs[10][62] ,
         \negative_inputs[10][61] , \negative_inputs[10][60] ,
         \negative_inputs[10][59] , \negative_inputs[10][58] ,
         \negative_inputs[10][57] , \negative_inputs[10][56] ,
         \negative_inputs[10][55] , \negative_inputs[10][54] ,
         \negative_inputs[10][53] , \negative_inputs[10][52] ,
         \negative_inputs[10][51] , \negative_inputs[10][50] ,
         \negative_inputs[10][49] , \negative_inputs[10][48] ,
         \negative_inputs[10][47] , \negative_inputs[10][46] ,
         \negative_inputs[10][45] , \negative_inputs[10][44] ,
         \negative_inputs[10][43] , \negative_inputs[10][42] ,
         \negative_inputs[10][41] , \negative_inputs[10][40] ,
         \negative_inputs[10][39] , \negative_inputs[10][38] ,
         \negative_inputs[10][37] , \negative_inputs[10][36] ,
         \negative_inputs[10][35] , \negative_inputs[10][34] ,
         \negative_inputs[10][33] , \negative_inputs[10][32] ,
         \negative_inputs[10][31] , \negative_inputs[10][30] ,
         \negative_inputs[10][29] , \negative_inputs[10][28] ,
         \negative_inputs[10][27] , \negative_inputs[10][26] ,
         \negative_inputs[10][25] , \negative_inputs[10][24] ,
         \negative_inputs[10][23] , \negative_inputs[10][22] ,
         \negative_inputs[10][21] , \negative_inputs[10][20] ,
         \negative_inputs[10][19] , \negative_inputs[10][18] ,
         \negative_inputs[10][17] , \negative_inputs[10][16] ,
         \negative_inputs[10][15] , \negative_inputs[10][14] ,
         \negative_inputs[10][13] , \negative_inputs[10][12] ,
         \negative_inputs[10][11] , \negative_inputs[10][10] ,
         \negative_inputs[10][9] , \negative_inputs[10][8] ,
         \negative_inputs[10][7] , \negative_inputs[10][6] ,
         \negative_inputs[10][5] , \negative_inputs[10][4] ,
         \negative_inputs[10][3] , \negative_inputs[10][2] ,
         \negative_inputs[10][1] , \negative_inputs[10][0] ,
         \negative_inputs[9][63] , \negative_inputs[9][62] ,
         \negative_inputs[9][61] , \negative_inputs[9][60] ,
         \negative_inputs[9][59] , \negative_inputs[9][58] ,
         \negative_inputs[9][57] , \negative_inputs[9][56] ,
         \negative_inputs[9][55] , \negative_inputs[9][54] ,
         \negative_inputs[9][53] , \negative_inputs[9][52] ,
         \negative_inputs[9][51] , \negative_inputs[9][50] ,
         \negative_inputs[9][49] , \negative_inputs[9][48] ,
         \negative_inputs[9][47] , \negative_inputs[9][46] ,
         \negative_inputs[9][45] , \negative_inputs[9][44] ,
         \negative_inputs[9][43] , \negative_inputs[9][42] ,
         \negative_inputs[9][41] , \negative_inputs[9][40] ,
         \negative_inputs[9][39] , \negative_inputs[9][38] ,
         \negative_inputs[9][37] , \negative_inputs[9][36] ,
         \negative_inputs[9][35] , \negative_inputs[9][34] ,
         \negative_inputs[9][33] , \negative_inputs[9][32] ,
         \negative_inputs[9][31] , \negative_inputs[9][30] ,
         \negative_inputs[9][29] , \negative_inputs[9][28] ,
         \negative_inputs[9][27] , \negative_inputs[9][26] ,
         \negative_inputs[9][25] , \negative_inputs[9][24] ,
         \negative_inputs[9][23] , \negative_inputs[9][22] ,
         \negative_inputs[9][21] , \negative_inputs[9][20] ,
         \negative_inputs[9][19] , \negative_inputs[9][18] ,
         \negative_inputs[9][17] , \negative_inputs[9][16] ,
         \negative_inputs[9][15] , \negative_inputs[9][14] ,
         \negative_inputs[9][13] , \negative_inputs[9][12] ,
         \negative_inputs[9][11] , \negative_inputs[9][10] ,
         \negative_inputs[9][9] , \negative_inputs[9][8] ,
         \negative_inputs[9][7] , \negative_inputs[9][6] ,
         \negative_inputs[9][5] , \negative_inputs[9][4] ,
         \negative_inputs[9][3] , \negative_inputs[9][2] ,
         \negative_inputs[9][1] , \negative_inputs[9][0] ,
         \negative_inputs[8][63] , \negative_inputs[8][62] ,
         \negative_inputs[8][61] , \negative_inputs[8][60] ,
         \negative_inputs[8][59] , \negative_inputs[8][58] ,
         \negative_inputs[8][57] , \negative_inputs[8][56] ,
         \negative_inputs[8][55] , \negative_inputs[8][54] ,
         \negative_inputs[8][53] , \negative_inputs[8][52] ,
         \negative_inputs[8][51] , \negative_inputs[8][50] ,
         \negative_inputs[8][49] , \negative_inputs[8][48] ,
         \negative_inputs[8][47] , \negative_inputs[8][46] ,
         \negative_inputs[8][45] , \negative_inputs[8][44] ,
         \negative_inputs[8][43] , \negative_inputs[8][42] ,
         \negative_inputs[8][41] , \negative_inputs[8][40] ,
         \negative_inputs[8][39] , \negative_inputs[8][38] ,
         \negative_inputs[8][37] , \negative_inputs[8][36] ,
         \negative_inputs[8][35] , \negative_inputs[8][34] ,
         \negative_inputs[8][33] , \negative_inputs[8][32] ,
         \negative_inputs[8][31] , \negative_inputs[8][30] ,
         \negative_inputs[8][29] , \negative_inputs[8][28] ,
         \negative_inputs[8][27] , \negative_inputs[8][26] ,
         \negative_inputs[8][25] , \negative_inputs[8][24] ,
         \negative_inputs[8][23] , \negative_inputs[8][22] ,
         \negative_inputs[8][21] , \negative_inputs[8][20] ,
         \negative_inputs[8][19] , \negative_inputs[8][18] ,
         \negative_inputs[8][17] , \negative_inputs[8][16] ,
         \negative_inputs[8][15] , \negative_inputs[8][14] ,
         \negative_inputs[8][13] , \negative_inputs[8][12] ,
         \negative_inputs[8][11] , \negative_inputs[8][10] ,
         \negative_inputs[8][9] , \negative_inputs[8][8] ,
         \negative_inputs[8][7] , \negative_inputs[8][6] ,
         \negative_inputs[8][5] , \negative_inputs[8][4] ,
         \negative_inputs[8][3] , \negative_inputs[8][2] ,
         \negative_inputs[8][1] , \negative_inputs[8][0] ,
         \negative_inputs[7][63] , \negative_inputs[7][62] ,
         \negative_inputs[7][61] , \negative_inputs[7][60] ,
         \negative_inputs[7][59] , \negative_inputs[7][58] ,
         \negative_inputs[7][57] , \negative_inputs[7][56] ,
         \negative_inputs[7][55] , \negative_inputs[7][54] ,
         \negative_inputs[7][53] , \negative_inputs[7][52] ,
         \negative_inputs[7][51] , \negative_inputs[7][50] ,
         \negative_inputs[7][49] , \negative_inputs[7][48] ,
         \negative_inputs[7][47] , \negative_inputs[7][46] ,
         \negative_inputs[7][45] , \negative_inputs[7][44] ,
         \negative_inputs[7][43] , \negative_inputs[7][42] ,
         \negative_inputs[7][41] , \negative_inputs[7][40] ,
         \negative_inputs[7][39] , \negative_inputs[7][38] ,
         \negative_inputs[7][37] , \negative_inputs[7][36] ,
         \negative_inputs[7][35] , \negative_inputs[7][34] ,
         \negative_inputs[7][33] , \negative_inputs[7][32] ,
         \negative_inputs[7][31] , \negative_inputs[7][30] ,
         \negative_inputs[7][29] , \negative_inputs[7][28] ,
         \negative_inputs[7][27] , \negative_inputs[7][26] ,
         \negative_inputs[7][25] , \negative_inputs[7][24] ,
         \negative_inputs[7][23] , \negative_inputs[7][22] ,
         \negative_inputs[7][21] , \negative_inputs[7][20] ,
         \negative_inputs[7][19] , \negative_inputs[7][18] ,
         \negative_inputs[7][17] , \negative_inputs[7][16] ,
         \negative_inputs[7][15] , \negative_inputs[7][14] ,
         \negative_inputs[7][13] , \negative_inputs[7][12] ,
         \negative_inputs[7][11] , \negative_inputs[7][10] ,
         \negative_inputs[7][9] , \negative_inputs[7][8] ,
         \negative_inputs[7][7] , \negative_inputs[7][6] ,
         \negative_inputs[7][5] , \negative_inputs[7][4] ,
         \negative_inputs[7][3] , \negative_inputs[7][2] ,
         \negative_inputs[7][1] , \negative_inputs[7][0] ,
         \negative_inputs[6][63] , \negative_inputs[6][62] ,
         \negative_inputs[6][61] , \negative_inputs[6][60] ,
         \negative_inputs[6][59] , \negative_inputs[6][58] ,
         \negative_inputs[6][57] , \negative_inputs[6][56] ,
         \negative_inputs[6][55] , \negative_inputs[6][54] ,
         \negative_inputs[6][53] , \negative_inputs[6][52] ,
         \negative_inputs[6][51] , \negative_inputs[6][50] ,
         \negative_inputs[6][49] , \negative_inputs[6][48] ,
         \negative_inputs[6][47] , \negative_inputs[6][46] ,
         \negative_inputs[6][45] , \negative_inputs[6][44] ,
         \negative_inputs[6][43] , \negative_inputs[6][42] ,
         \negative_inputs[6][41] , \negative_inputs[6][40] ,
         \negative_inputs[6][39] , \negative_inputs[6][38] ,
         \negative_inputs[6][37] , \negative_inputs[6][36] ,
         \negative_inputs[6][35] , \negative_inputs[6][34] ,
         \negative_inputs[6][33] , \negative_inputs[6][32] ,
         \negative_inputs[6][31] , \negative_inputs[6][30] ,
         \negative_inputs[6][29] , \negative_inputs[6][28] ,
         \negative_inputs[6][27] , \negative_inputs[6][26] ,
         \negative_inputs[6][25] , \negative_inputs[6][24] ,
         \negative_inputs[6][23] , \negative_inputs[6][22] ,
         \negative_inputs[6][21] , \negative_inputs[6][20] ,
         \negative_inputs[6][19] , \negative_inputs[6][18] ,
         \negative_inputs[6][17] , \negative_inputs[6][16] ,
         \negative_inputs[6][15] , \negative_inputs[6][14] ,
         \negative_inputs[6][13] , \negative_inputs[6][12] ,
         \negative_inputs[6][11] , \negative_inputs[6][10] ,
         \negative_inputs[6][9] , \negative_inputs[6][8] ,
         \negative_inputs[6][7] , \negative_inputs[6][6] ,
         \negative_inputs[6][5] , \negative_inputs[6][4] ,
         \negative_inputs[6][3] , \negative_inputs[6][2] ,
         \negative_inputs[6][1] , \negative_inputs[6][0] ,
         \negative_inputs[5][63] , \negative_inputs[5][62] ,
         \negative_inputs[5][61] , \negative_inputs[5][60] ,
         \negative_inputs[5][59] , \negative_inputs[5][58] ,
         \negative_inputs[5][57] , \negative_inputs[5][56] ,
         \negative_inputs[5][55] , \negative_inputs[5][54] ,
         \negative_inputs[5][53] , \negative_inputs[5][52] ,
         \negative_inputs[5][51] , \negative_inputs[5][50] ,
         \negative_inputs[5][49] , \negative_inputs[5][48] ,
         \negative_inputs[5][47] , \negative_inputs[5][46] ,
         \negative_inputs[5][45] , \negative_inputs[5][44] ,
         \negative_inputs[5][43] , \negative_inputs[5][42] ,
         \negative_inputs[5][41] , \negative_inputs[5][40] ,
         \negative_inputs[5][39] , \negative_inputs[5][38] ,
         \negative_inputs[5][37] , \negative_inputs[5][36] ,
         \negative_inputs[5][35] , \negative_inputs[5][34] ,
         \negative_inputs[5][33] , \negative_inputs[5][32] ,
         \negative_inputs[5][31] , \negative_inputs[5][30] ,
         \negative_inputs[5][29] , \negative_inputs[5][28] ,
         \negative_inputs[5][27] , \negative_inputs[5][26] ,
         \negative_inputs[5][25] , \negative_inputs[5][24] ,
         \negative_inputs[5][23] , \negative_inputs[5][22] ,
         \negative_inputs[5][21] , \negative_inputs[5][20] ,
         \negative_inputs[5][19] , \negative_inputs[5][18] ,
         \negative_inputs[5][17] , \negative_inputs[5][16] ,
         \negative_inputs[5][15] , \negative_inputs[5][14] ,
         \negative_inputs[5][13] , \negative_inputs[5][12] ,
         \negative_inputs[5][11] , \negative_inputs[5][10] ,
         \negative_inputs[5][9] , \negative_inputs[5][8] ,
         \negative_inputs[5][7] , \negative_inputs[5][6] ,
         \negative_inputs[5][5] , \negative_inputs[5][4] ,
         \negative_inputs[5][3] , \negative_inputs[5][2] ,
         \negative_inputs[5][1] , \negative_inputs[5][0] ,
         \negative_inputs[4][63] , \negative_inputs[4][62] ,
         \negative_inputs[4][61] , \negative_inputs[4][60] ,
         \negative_inputs[4][59] , \negative_inputs[4][58] ,
         \negative_inputs[4][57] , \negative_inputs[4][56] ,
         \negative_inputs[4][55] , \negative_inputs[4][54] ,
         \negative_inputs[4][53] , \negative_inputs[4][52] ,
         \negative_inputs[4][51] , \negative_inputs[4][50] ,
         \negative_inputs[4][49] , \negative_inputs[4][48] ,
         \negative_inputs[4][47] , \negative_inputs[4][46] ,
         \negative_inputs[4][45] , \negative_inputs[4][44] ,
         \negative_inputs[4][43] , \negative_inputs[4][42] ,
         \negative_inputs[4][41] , \negative_inputs[4][40] ,
         \negative_inputs[4][39] , \negative_inputs[4][38] ,
         \negative_inputs[4][37] , \negative_inputs[4][36] ,
         \negative_inputs[4][35] , \negative_inputs[4][34] ,
         \negative_inputs[4][33] , \negative_inputs[4][32] ,
         \negative_inputs[4][31] , \negative_inputs[4][30] ,
         \negative_inputs[4][29] , \negative_inputs[4][28] ,
         \negative_inputs[4][27] , \negative_inputs[4][26] ,
         \negative_inputs[4][25] , \negative_inputs[4][24] ,
         \negative_inputs[4][23] , \negative_inputs[4][22] ,
         \negative_inputs[4][21] , \negative_inputs[4][20] ,
         \negative_inputs[4][19] , \negative_inputs[4][18] ,
         \negative_inputs[4][17] , \negative_inputs[4][16] ,
         \negative_inputs[4][15] , \negative_inputs[4][14] ,
         \negative_inputs[4][13] , \negative_inputs[4][12] ,
         \negative_inputs[4][11] , \negative_inputs[4][10] ,
         \negative_inputs[4][9] , \negative_inputs[4][8] ,
         \negative_inputs[4][7] , \negative_inputs[4][6] ,
         \negative_inputs[4][5] , \negative_inputs[4][4] ,
         \negative_inputs[4][3] , \negative_inputs[4][2] ,
         \negative_inputs[4][1] , \negative_inputs[4][0] ,
         \negative_inputs[3][63] , \negative_inputs[3][62] ,
         \negative_inputs[3][61] , \negative_inputs[3][60] ,
         \negative_inputs[3][59] , \negative_inputs[3][58] ,
         \negative_inputs[3][57] , \negative_inputs[3][56] ,
         \negative_inputs[3][55] , \negative_inputs[3][54] ,
         \negative_inputs[3][53] , \negative_inputs[3][52] ,
         \negative_inputs[3][51] , \negative_inputs[3][50] ,
         \negative_inputs[3][49] , \negative_inputs[3][48] ,
         \negative_inputs[3][47] , \negative_inputs[3][46] ,
         \negative_inputs[3][45] , \negative_inputs[3][44] ,
         \negative_inputs[3][43] , \negative_inputs[3][42] ,
         \negative_inputs[3][41] , \negative_inputs[3][40] ,
         \negative_inputs[3][39] , \negative_inputs[3][38] ,
         \negative_inputs[3][37] , \negative_inputs[3][36] ,
         \negative_inputs[3][35] , \negative_inputs[3][34] ,
         \negative_inputs[3][33] , \negative_inputs[3][32] ,
         \negative_inputs[3][31] , \negative_inputs[3][30] ,
         \negative_inputs[3][29] , \negative_inputs[3][28] ,
         \negative_inputs[3][27] , \negative_inputs[3][26] ,
         \negative_inputs[3][25] , \negative_inputs[3][24] ,
         \negative_inputs[3][23] , \negative_inputs[3][22] ,
         \negative_inputs[3][21] , \negative_inputs[3][20] ,
         \negative_inputs[3][19] , \negative_inputs[3][18] ,
         \negative_inputs[3][17] , \negative_inputs[3][16] ,
         \negative_inputs[3][15] , \negative_inputs[3][14] ,
         \negative_inputs[3][13] , \negative_inputs[3][12] ,
         \negative_inputs[3][11] , \negative_inputs[3][10] ,
         \negative_inputs[3][9] , \negative_inputs[3][8] ,
         \negative_inputs[3][7] , \negative_inputs[3][6] ,
         \negative_inputs[3][5] , \negative_inputs[3][4] ,
         \negative_inputs[3][3] , \negative_inputs[3][2] ,
         \negative_inputs[3][1] , \negative_inputs[3][0] ,
         \negative_inputs[2][63] , \negative_inputs[2][62] ,
         \negative_inputs[2][61] , \negative_inputs[2][60] ,
         \negative_inputs[2][59] , \negative_inputs[2][58] ,
         \negative_inputs[2][57] , \negative_inputs[2][56] ,
         \negative_inputs[2][55] , \negative_inputs[2][54] ,
         \negative_inputs[2][53] , \negative_inputs[2][52] ,
         \negative_inputs[2][51] , \negative_inputs[2][50] ,
         \negative_inputs[2][49] , \negative_inputs[2][48] ,
         \negative_inputs[2][47] , \negative_inputs[2][46] ,
         \negative_inputs[2][45] , \negative_inputs[2][44] ,
         \negative_inputs[2][43] , \negative_inputs[2][42] ,
         \negative_inputs[2][41] , \negative_inputs[2][40] ,
         \negative_inputs[2][39] , \negative_inputs[2][38] ,
         \negative_inputs[2][37] , \negative_inputs[2][36] ,
         \negative_inputs[2][35] , \negative_inputs[2][34] ,
         \negative_inputs[2][33] , \negative_inputs[2][32] ,
         \negative_inputs[2][31] , \negative_inputs[2][30] ,
         \negative_inputs[2][29] , \negative_inputs[2][28] ,
         \negative_inputs[2][27] , \negative_inputs[2][26] ,
         \negative_inputs[2][25] , \negative_inputs[2][24] ,
         \negative_inputs[2][23] , \negative_inputs[2][22] ,
         \negative_inputs[2][21] , \negative_inputs[2][20] ,
         \negative_inputs[2][19] , \negative_inputs[2][18] ,
         \negative_inputs[2][17] , \negative_inputs[2][16] ,
         \negative_inputs[2][15] , \negative_inputs[2][14] ,
         \negative_inputs[2][13] , \negative_inputs[2][12] ,
         \negative_inputs[2][11] , \negative_inputs[2][10] ,
         \negative_inputs[2][9] , \negative_inputs[2][8] ,
         \negative_inputs[2][7] , \negative_inputs[2][6] ,
         \negative_inputs[2][5] , \negative_inputs[2][4] ,
         \negative_inputs[2][3] , \negative_inputs[2][2] ,
         \negative_inputs[2][1] , \negative_inputs[2][0] ,
         \negative_inputs[1][63] , \negative_inputs[1][62] ,
         \negative_inputs[1][61] , \negative_inputs[1][60] ,
         \negative_inputs[1][59] , \negative_inputs[1][58] ,
         \negative_inputs[1][57] , \negative_inputs[1][56] ,
         \negative_inputs[1][55] , \negative_inputs[1][54] ,
         \negative_inputs[1][53] , \negative_inputs[1][52] ,
         \negative_inputs[1][51] , \negative_inputs[1][50] ,
         \negative_inputs[1][49] , \negative_inputs[1][48] ,
         \negative_inputs[1][47] , \negative_inputs[1][46] ,
         \negative_inputs[1][45] , \negative_inputs[1][44] ,
         \negative_inputs[1][43] , \negative_inputs[1][42] ,
         \negative_inputs[1][41] , \negative_inputs[1][40] ,
         \negative_inputs[1][39] , \negative_inputs[1][38] ,
         \negative_inputs[1][37] , \negative_inputs[1][36] ,
         \negative_inputs[1][35] , \negative_inputs[1][34] ,
         \negative_inputs[1][33] , \negative_inputs[1][32] ,
         \negative_inputs[1][31] , \negative_inputs[1][30] ,
         \negative_inputs[1][29] , \negative_inputs[1][28] ,
         \negative_inputs[1][27] , \negative_inputs[1][26] ,
         \negative_inputs[1][25] , \negative_inputs[1][24] ,
         \negative_inputs[1][23] , \negative_inputs[1][22] ,
         \negative_inputs[1][21] , \negative_inputs[1][20] ,
         \negative_inputs[1][19] , \negative_inputs[1][18] ,
         \negative_inputs[1][17] , \negative_inputs[1][16] ,
         \negative_inputs[1][15] , \negative_inputs[1][14] ,
         \negative_inputs[1][13] , \negative_inputs[1][12] ,
         \negative_inputs[1][11] , \negative_inputs[1][10] ,
         \negative_inputs[1][9] , \negative_inputs[1][8] ,
         \negative_inputs[1][7] , \negative_inputs[1][6] ,
         \negative_inputs[1][5] , \negative_inputs[1][4] ,
         \negative_inputs[1][3] , \negative_inputs[1][2] ,
         \negative_inputs[1][1] , \negative_inputs[1][0] ,
         \negative_inputs[0][63] , \negative_inputs[0][62] ,
         \negative_inputs[0][61] , \negative_inputs[0][60] ,
         \negative_inputs[0][59] , \negative_inputs[0][58] ,
         \negative_inputs[0][57] , \negative_inputs[0][56] ,
         \negative_inputs[0][55] , \negative_inputs[0][54] ,
         \negative_inputs[0][53] , \negative_inputs[0][52] ,
         \negative_inputs[0][51] , \negative_inputs[0][50] ,
         \negative_inputs[0][49] , \negative_inputs[0][48] ,
         \negative_inputs[0][47] , \negative_inputs[0][46] ,
         \negative_inputs[0][45] , \negative_inputs[0][44] ,
         \negative_inputs[0][43] , \negative_inputs[0][42] ,
         \negative_inputs[0][41] , \negative_inputs[0][40] ,
         \negative_inputs[0][39] , \negative_inputs[0][38] ,
         \negative_inputs[0][37] , \negative_inputs[0][36] ,
         \negative_inputs[0][35] , \negative_inputs[0][34] ,
         \negative_inputs[0][33] , \negative_inputs[0][32] ,
         \negative_inputs[0][31] , \negative_inputs[0][30] ,
         \negative_inputs[0][29] , \negative_inputs[0][28] ,
         \negative_inputs[0][27] , \negative_inputs[0][26] ,
         \negative_inputs[0][25] , \negative_inputs[0][24] ,
         \negative_inputs[0][23] , \negative_inputs[0][22] ,
         \negative_inputs[0][21] , \negative_inputs[0][20] ,
         \negative_inputs[0][19] , \negative_inputs[0][18] ,
         \negative_inputs[0][17] , \negative_inputs[0][16] ,
         \negative_inputs[0][15] , \negative_inputs[0][14] ,
         \negative_inputs[0][13] , \negative_inputs[0][12] ,
         \negative_inputs[0][11] , \negative_inputs[0][10] ,
         \negative_inputs[0][9] , \negative_inputs[0][8] ,
         \negative_inputs[0][7] , \negative_inputs[0][6] ,
         \negative_inputs[0][5] , \negative_inputs[0][4] ,
         \negative_inputs[0][3] , \negative_inputs[0][2] ,
         \negative_inputs[0][1] , \negative_inputs[0][0] ,
         \ADDER_IN_from_mux[15][63] , \ADDER_IN_from_mux[15][62] ,
         \ADDER_IN_from_mux[15][61] , \ADDER_IN_from_mux[15][60] ,
         \ADDER_IN_from_mux[15][59] , \ADDER_IN_from_mux[15][58] ,
         \ADDER_IN_from_mux[15][57] , \ADDER_IN_from_mux[15][56] ,
         \ADDER_IN_from_mux[15][55] , \ADDER_IN_from_mux[15][54] ,
         \ADDER_IN_from_mux[15][53] , \ADDER_IN_from_mux[15][52] ,
         \ADDER_IN_from_mux[15][51] , \ADDER_IN_from_mux[15][50] ,
         \ADDER_IN_from_mux[15][49] , \ADDER_IN_from_mux[15][48] ,
         \ADDER_IN_from_mux[15][47] , \ADDER_IN_from_mux[15][46] ,
         \ADDER_IN_from_mux[15][45] , \ADDER_IN_from_mux[15][44] ,
         \ADDER_IN_from_mux[15][43] , \ADDER_IN_from_mux[15][42] ,
         \ADDER_IN_from_mux[15][41] , \ADDER_IN_from_mux[15][40] ,
         \ADDER_IN_from_mux[15][39] , \ADDER_IN_from_mux[15][38] ,
         \ADDER_IN_from_mux[15][37] , \ADDER_IN_from_mux[15][36] ,
         \ADDER_IN_from_mux[15][35] , \ADDER_IN_from_mux[15][34] ,
         \ADDER_IN_from_mux[15][33] , \ADDER_IN_from_mux[15][32] ,
         \ADDER_IN_from_mux[15][31] , \ADDER_IN_from_mux[15][30] ,
         \ADDER_IN_from_mux[15][29] , \ADDER_IN_from_mux[15][28] ,
         \ADDER_IN_from_mux[15][27] , \ADDER_IN_from_mux[15][26] ,
         \ADDER_IN_from_mux[15][25] , \ADDER_IN_from_mux[15][24] ,
         \ADDER_IN_from_mux[15][23] , \ADDER_IN_from_mux[15][22] ,
         \ADDER_IN_from_mux[15][21] , \ADDER_IN_from_mux[15][20] ,
         \ADDER_IN_from_mux[15][19] , \ADDER_IN_from_mux[15][18] ,
         \ADDER_IN_from_mux[15][17] , \ADDER_IN_from_mux[15][16] ,
         \ADDER_IN_from_mux[15][15] , \ADDER_IN_from_mux[15][14] ,
         \ADDER_IN_from_mux[15][13] , \ADDER_IN_from_mux[15][12] ,
         \ADDER_IN_from_mux[15][11] , \ADDER_IN_from_mux[15][10] ,
         \ADDER_IN_from_mux[15][9] , \ADDER_IN_from_mux[15][8] ,
         \ADDER_IN_from_mux[15][7] , \ADDER_IN_from_mux[15][6] ,
         \ADDER_IN_from_mux[15][5] , \ADDER_IN_from_mux[15][4] ,
         \ADDER_IN_from_mux[15][3] , \ADDER_IN_from_mux[15][2] ,
         \ADDER_IN_from_mux[15][1] , \ADDER_IN_from_mux[15][0] ,
         \ADDER_IN_from_mux[14][63] , \ADDER_IN_from_mux[14][62] ,
         \ADDER_IN_from_mux[14][61] , \ADDER_IN_from_mux[14][60] ,
         \ADDER_IN_from_mux[14][59] , \ADDER_IN_from_mux[14][58] ,
         \ADDER_IN_from_mux[14][57] , \ADDER_IN_from_mux[14][56] ,
         \ADDER_IN_from_mux[14][55] , \ADDER_IN_from_mux[14][54] ,
         \ADDER_IN_from_mux[14][53] , \ADDER_IN_from_mux[14][52] ,
         \ADDER_IN_from_mux[14][51] , \ADDER_IN_from_mux[14][50] ,
         \ADDER_IN_from_mux[14][49] , \ADDER_IN_from_mux[14][48] ,
         \ADDER_IN_from_mux[14][47] , \ADDER_IN_from_mux[14][46] ,
         \ADDER_IN_from_mux[14][45] , \ADDER_IN_from_mux[14][44] ,
         \ADDER_IN_from_mux[14][43] , \ADDER_IN_from_mux[14][42] ,
         \ADDER_IN_from_mux[14][41] , \ADDER_IN_from_mux[14][40] ,
         \ADDER_IN_from_mux[14][39] , \ADDER_IN_from_mux[14][38] ,
         \ADDER_IN_from_mux[14][37] , \ADDER_IN_from_mux[14][36] ,
         \ADDER_IN_from_mux[14][35] , \ADDER_IN_from_mux[14][34] ,
         \ADDER_IN_from_mux[14][33] , \ADDER_IN_from_mux[14][32] ,
         \ADDER_IN_from_mux[14][31] , \ADDER_IN_from_mux[14][30] ,
         \ADDER_IN_from_mux[14][29] , \ADDER_IN_from_mux[14][28] ,
         \ADDER_IN_from_mux[14][27] , \ADDER_IN_from_mux[14][26] ,
         \ADDER_IN_from_mux[14][25] , \ADDER_IN_from_mux[14][24] ,
         \ADDER_IN_from_mux[14][23] , \ADDER_IN_from_mux[14][22] ,
         \ADDER_IN_from_mux[14][21] , \ADDER_IN_from_mux[14][20] ,
         \ADDER_IN_from_mux[14][19] , \ADDER_IN_from_mux[14][18] ,
         \ADDER_IN_from_mux[14][17] , \ADDER_IN_from_mux[14][16] ,
         \ADDER_IN_from_mux[14][15] , \ADDER_IN_from_mux[14][14] ,
         \ADDER_IN_from_mux[14][13] , \ADDER_IN_from_mux[14][12] ,
         \ADDER_IN_from_mux[14][11] , \ADDER_IN_from_mux[14][10] ,
         \ADDER_IN_from_mux[14][9] , \ADDER_IN_from_mux[14][8] ,
         \ADDER_IN_from_mux[14][7] , \ADDER_IN_from_mux[14][6] ,
         \ADDER_IN_from_mux[14][5] , \ADDER_IN_from_mux[14][4] ,
         \ADDER_IN_from_mux[14][3] , \ADDER_IN_from_mux[14][2] ,
         \ADDER_IN_from_mux[14][1] , \ADDER_IN_from_mux[14][0] ,
         \ADDER_IN_from_mux[13][63] , \ADDER_IN_from_mux[13][62] ,
         \ADDER_IN_from_mux[13][61] , \ADDER_IN_from_mux[13][60] ,
         \ADDER_IN_from_mux[13][59] , \ADDER_IN_from_mux[13][58] ,
         \ADDER_IN_from_mux[13][57] , \ADDER_IN_from_mux[13][56] ,
         \ADDER_IN_from_mux[13][55] , \ADDER_IN_from_mux[13][54] ,
         \ADDER_IN_from_mux[13][53] , \ADDER_IN_from_mux[13][52] ,
         \ADDER_IN_from_mux[13][51] , \ADDER_IN_from_mux[13][50] ,
         \ADDER_IN_from_mux[13][49] , \ADDER_IN_from_mux[13][48] ,
         \ADDER_IN_from_mux[13][47] , \ADDER_IN_from_mux[13][46] ,
         \ADDER_IN_from_mux[13][45] , \ADDER_IN_from_mux[13][44] ,
         \ADDER_IN_from_mux[13][43] , \ADDER_IN_from_mux[13][42] ,
         \ADDER_IN_from_mux[13][41] , \ADDER_IN_from_mux[13][40] ,
         \ADDER_IN_from_mux[13][39] , \ADDER_IN_from_mux[13][38] ,
         \ADDER_IN_from_mux[13][37] , \ADDER_IN_from_mux[13][36] ,
         \ADDER_IN_from_mux[13][35] , \ADDER_IN_from_mux[13][34] ,
         \ADDER_IN_from_mux[13][33] , \ADDER_IN_from_mux[13][32] ,
         \ADDER_IN_from_mux[13][31] , \ADDER_IN_from_mux[13][30] ,
         \ADDER_IN_from_mux[13][29] , \ADDER_IN_from_mux[13][28] ,
         \ADDER_IN_from_mux[13][27] , \ADDER_IN_from_mux[13][26] ,
         \ADDER_IN_from_mux[13][25] , \ADDER_IN_from_mux[13][24] ,
         \ADDER_IN_from_mux[13][23] , \ADDER_IN_from_mux[13][22] ,
         \ADDER_IN_from_mux[13][21] , \ADDER_IN_from_mux[13][20] ,
         \ADDER_IN_from_mux[13][19] , \ADDER_IN_from_mux[13][18] ,
         \ADDER_IN_from_mux[13][17] , \ADDER_IN_from_mux[13][16] ,
         \ADDER_IN_from_mux[13][15] , \ADDER_IN_from_mux[13][14] ,
         \ADDER_IN_from_mux[13][13] , \ADDER_IN_from_mux[13][12] ,
         \ADDER_IN_from_mux[13][11] , \ADDER_IN_from_mux[13][10] ,
         \ADDER_IN_from_mux[13][9] , \ADDER_IN_from_mux[13][8] ,
         \ADDER_IN_from_mux[13][7] , \ADDER_IN_from_mux[13][6] ,
         \ADDER_IN_from_mux[13][5] , \ADDER_IN_from_mux[13][4] ,
         \ADDER_IN_from_mux[13][3] , \ADDER_IN_from_mux[13][2] ,
         \ADDER_IN_from_mux[13][1] , \ADDER_IN_from_mux[13][0] ,
         \ADDER_IN_from_mux[12][63] , \ADDER_IN_from_mux[12][62] ,
         \ADDER_IN_from_mux[12][61] , \ADDER_IN_from_mux[12][60] ,
         \ADDER_IN_from_mux[12][59] , \ADDER_IN_from_mux[12][58] ,
         \ADDER_IN_from_mux[12][57] , \ADDER_IN_from_mux[12][56] ,
         \ADDER_IN_from_mux[12][55] , \ADDER_IN_from_mux[12][54] ,
         \ADDER_IN_from_mux[12][53] , \ADDER_IN_from_mux[12][52] ,
         \ADDER_IN_from_mux[12][51] , \ADDER_IN_from_mux[12][50] ,
         \ADDER_IN_from_mux[12][49] , \ADDER_IN_from_mux[12][48] ,
         \ADDER_IN_from_mux[12][47] , \ADDER_IN_from_mux[12][46] ,
         \ADDER_IN_from_mux[12][45] , \ADDER_IN_from_mux[12][44] ,
         \ADDER_IN_from_mux[12][43] , \ADDER_IN_from_mux[12][42] ,
         \ADDER_IN_from_mux[12][41] , \ADDER_IN_from_mux[12][40] ,
         \ADDER_IN_from_mux[12][39] , \ADDER_IN_from_mux[12][38] ,
         \ADDER_IN_from_mux[12][37] , \ADDER_IN_from_mux[12][36] ,
         \ADDER_IN_from_mux[12][35] , \ADDER_IN_from_mux[12][34] ,
         \ADDER_IN_from_mux[12][33] , \ADDER_IN_from_mux[12][32] ,
         \ADDER_IN_from_mux[12][31] , \ADDER_IN_from_mux[12][30] ,
         \ADDER_IN_from_mux[12][29] , \ADDER_IN_from_mux[12][28] ,
         \ADDER_IN_from_mux[12][27] , \ADDER_IN_from_mux[12][26] ,
         \ADDER_IN_from_mux[12][25] , \ADDER_IN_from_mux[12][24] ,
         \ADDER_IN_from_mux[12][23] , \ADDER_IN_from_mux[12][22] ,
         \ADDER_IN_from_mux[12][21] , \ADDER_IN_from_mux[12][20] ,
         \ADDER_IN_from_mux[12][19] , \ADDER_IN_from_mux[12][18] ,
         \ADDER_IN_from_mux[12][17] , \ADDER_IN_from_mux[12][16] ,
         \ADDER_IN_from_mux[12][15] , \ADDER_IN_from_mux[12][14] ,
         \ADDER_IN_from_mux[12][13] , \ADDER_IN_from_mux[12][12] ,
         \ADDER_IN_from_mux[12][11] , \ADDER_IN_from_mux[12][10] ,
         \ADDER_IN_from_mux[12][9] , \ADDER_IN_from_mux[12][8] ,
         \ADDER_IN_from_mux[12][7] , \ADDER_IN_from_mux[12][6] ,
         \ADDER_IN_from_mux[12][5] , \ADDER_IN_from_mux[12][4] ,
         \ADDER_IN_from_mux[12][3] , \ADDER_IN_from_mux[12][2] ,
         \ADDER_IN_from_mux[12][1] , \ADDER_IN_from_mux[12][0] ,
         \ADDER_IN_from_mux[11][63] , \ADDER_IN_from_mux[11][62] ,
         \ADDER_IN_from_mux[11][61] , \ADDER_IN_from_mux[11][60] ,
         \ADDER_IN_from_mux[11][59] , \ADDER_IN_from_mux[11][58] ,
         \ADDER_IN_from_mux[11][57] , \ADDER_IN_from_mux[11][56] ,
         \ADDER_IN_from_mux[11][55] , \ADDER_IN_from_mux[11][54] ,
         \ADDER_IN_from_mux[11][53] , \ADDER_IN_from_mux[11][52] ,
         \ADDER_IN_from_mux[11][51] , \ADDER_IN_from_mux[11][50] ,
         \ADDER_IN_from_mux[11][49] , \ADDER_IN_from_mux[11][48] ,
         \ADDER_IN_from_mux[11][47] , \ADDER_IN_from_mux[11][46] ,
         \ADDER_IN_from_mux[11][45] , \ADDER_IN_from_mux[11][44] ,
         \ADDER_IN_from_mux[11][43] , \ADDER_IN_from_mux[11][42] ,
         \ADDER_IN_from_mux[11][41] , \ADDER_IN_from_mux[11][40] ,
         \ADDER_IN_from_mux[11][39] , \ADDER_IN_from_mux[11][38] ,
         \ADDER_IN_from_mux[11][37] , \ADDER_IN_from_mux[11][36] ,
         \ADDER_IN_from_mux[11][35] , \ADDER_IN_from_mux[11][34] ,
         \ADDER_IN_from_mux[11][33] , \ADDER_IN_from_mux[11][32] ,
         \ADDER_IN_from_mux[11][31] , \ADDER_IN_from_mux[11][30] ,
         \ADDER_IN_from_mux[11][29] , \ADDER_IN_from_mux[11][28] ,
         \ADDER_IN_from_mux[11][27] , \ADDER_IN_from_mux[11][26] ,
         \ADDER_IN_from_mux[11][25] , \ADDER_IN_from_mux[11][24] ,
         \ADDER_IN_from_mux[11][23] , \ADDER_IN_from_mux[11][22] ,
         \ADDER_IN_from_mux[11][21] , \ADDER_IN_from_mux[11][20] ,
         \ADDER_IN_from_mux[11][19] , \ADDER_IN_from_mux[11][18] ,
         \ADDER_IN_from_mux[11][17] , \ADDER_IN_from_mux[11][16] ,
         \ADDER_IN_from_mux[11][15] , \ADDER_IN_from_mux[11][14] ,
         \ADDER_IN_from_mux[11][13] , \ADDER_IN_from_mux[11][12] ,
         \ADDER_IN_from_mux[11][11] , \ADDER_IN_from_mux[11][10] ,
         \ADDER_IN_from_mux[11][9] , \ADDER_IN_from_mux[11][8] ,
         \ADDER_IN_from_mux[11][7] , \ADDER_IN_from_mux[11][6] ,
         \ADDER_IN_from_mux[11][5] , \ADDER_IN_from_mux[11][4] ,
         \ADDER_IN_from_mux[11][3] , \ADDER_IN_from_mux[11][2] ,
         \ADDER_IN_from_mux[11][1] , \ADDER_IN_from_mux[11][0] ,
         \ADDER_IN_from_mux[10][63] , \ADDER_IN_from_mux[10][62] ,
         \ADDER_IN_from_mux[10][61] , \ADDER_IN_from_mux[10][60] ,
         \ADDER_IN_from_mux[10][59] , \ADDER_IN_from_mux[10][58] ,
         \ADDER_IN_from_mux[10][57] , \ADDER_IN_from_mux[10][56] ,
         \ADDER_IN_from_mux[10][55] , \ADDER_IN_from_mux[10][54] ,
         \ADDER_IN_from_mux[10][53] , \ADDER_IN_from_mux[10][52] ,
         \ADDER_IN_from_mux[10][51] , \ADDER_IN_from_mux[10][50] ,
         \ADDER_IN_from_mux[10][49] , \ADDER_IN_from_mux[10][48] ,
         \ADDER_IN_from_mux[10][47] , \ADDER_IN_from_mux[10][46] ,
         \ADDER_IN_from_mux[10][45] , \ADDER_IN_from_mux[10][44] ,
         \ADDER_IN_from_mux[10][43] , \ADDER_IN_from_mux[10][42] ,
         \ADDER_IN_from_mux[10][41] , \ADDER_IN_from_mux[10][40] ,
         \ADDER_IN_from_mux[10][39] , \ADDER_IN_from_mux[10][38] ,
         \ADDER_IN_from_mux[10][37] , \ADDER_IN_from_mux[10][36] ,
         \ADDER_IN_from_mux[10][35] , \ADDER_IN_from_mux[10][34] ,
         \ADDER_IN_from_mux[10][33] , \ADDER_IN_from_mux[10][32] ,
         \ADDER_IN_from_mux[10][31] , \ADDER_IN_from_mux[10][30] ,
         \ADDER_IN_from_mux[10][29] , \ADDER_IN_from_mux[10][28] ,
         \ADDER_IN_from_mux[10][27] , \ADDER_IN_from_mux[10][26] ,
         \ADDER_IN_from_mux[10][25] , \ADDER_IN_from_mux[10][24] ,
         \ADDER_IN_from_mux[10][23] , \ADDER_IN_from_mux[10][22] ,
         \ADDER_IN_from_mux[10][21] , \ADDER_IN_from_mux[10][20] ,
         \ADDER_IN_from_mux[10][19] , \ADDER_IN_from_mux[10][18] ,
         \ADDER_IN_from_mux[10][17] , \ADDER_IN_from_mux[10][16] ,
         \ADDER_IN_from_mux[10][15] , \ADDER_IN_from_mux[10][14] ,
         \ADDER_IN_from_mux[10][13] , \ADDER_IN_from_mux[10][12] ,
         \ADDER_IN_from_mux[10][11] , \ADDER_IN_from_mux[10][10] ,
         \ADDER_IN_from_mux[10][9] , \ADDER_IN_from_mux[10][8] ,
         \ADDER_IN_from_mux[10][7] , \ADDER_IN_from_mux[10][6] ,
         \ADDER_IN_from_mux[10][5] , \ADDER_IN_from_mux[10][4] ,
         \ADDER_IN_from_mux[10][3] , \ADDER_IN_from_mux[10][2] ,
         \ADDER_IN_from_mux[10][1] , \ADDER_IN_from_mux[10][0] ,
         \ADDER_IN_from_mux[9][63] , \ADDER_IN_from_mux[9][62] ,
         \ADDER_IN_from_mux[9][61] , \ADDER_IN_from_mux[9][60] ,
         \ADDER_IN_from_mux[9][59] , \ADDER_IN_from_mux[9][58] ,
         \ADDER_IN_from_mux[9][57] , \ADDER_IN_from_mux[9][56] ,
         \ADDER_IN_from_mux[9][55] , \ADDER_IN_from_mux[9][54] ,
         \ADDER_IN_from_mux[9][53] , \ADDER_IN_from_mux[9][52] ,
         \ADDER_IN_from_mux[9][51] , \ADDER_IN_from_mux[9][50] ,
         \ADDER_IN_from_mux[9][49] , \ADDER_IN_from_mux[9][48] ,
         \ADDER_IN_from_mux[9][47] , \ADDER_IN_from_mux[9][46] ,
         \ADDER_IN_from_mux[9][45] , \ADDER_IN_from_mux[9][44] ,
         \ADDER_IN_from_mux[9][43] , \ADDER_IN_from_mux[9][42] ,
         \ADDER_IN_from_mux[9][41] , \ADDER_IN_from_mux[9][40] ,
         \ADDER_IN_from_mux[9][39] , \ADDER_IN_from_mux[9][38] ,
         \ADDER_IN_from_mux[9][37] , \ADDER_IN_from_mux[9][36] ,
         \ADDER_IN_from_mux[9][35] , \ADDER_IN_from_mux[9][34] ,
         \ADDER_IN_from_mux[9][33] , \ADDER_IN_from_mux[9][32] ,
         \ADDER_IN_from_mux[9][31] , \ADDER_IN_from_mux[9][30] ,
         \ADDER_IN_from_mux[9][29] , \ADDER_IN_from_mux[9][28] ,
         \ADDER_IN_from_mux[9][27] , \ADDER_IN_from_mux[9][26] ,
         \ADDER_IN_from_mux[9][25] , \ADDER_IN_from_mux[9][24] ,
         \ADDER_IN_from_mux[9][23] , \ADDER_IN_from_mux[9][22] ,
         \ADDER_IN_from_mux[9][21] , \ADDER_IN_from_mux[9][20] ,
         \ADDER_IN_from_mux[9][19] , \ADDER_IN_from_mux[9][18] ,
         \ADDER_IN_from_mux[9][17] , \ADDER_IN_from_mux[9][16] ,
         \ADDER_IN_from_mux[9][15] , \ADDER_IN_from_mux[9][14] ,
         \ADDER_IN_from_mux[9][13] , \ADDER_IN_from_mux[9][12] ,
         \ADDER_IN_from_mux[9][11] , \ADDER_IN_from_mux[9][10] ,
         \ADDER_IN_from_mux[9][9] , \ADDER_IN_from_mux[9][8] ,
         \ADDER_IN_from_mux[9][7] , \ADDER_IN_from_mux[9][6] ,
         \ADDER_IN_from_mux[9][5] , \ADDER_IN_from_mux[9][4] ,
         \ADDER_IN_from_mux[9][3] , \ADDER_IN_from_mux[9][2] ,
         \ADDER_IN_from_mux[9][1] , \ADDER_IN_from_mux[9][0] ,
         \ADDER_IN_from_mux[8][63] , \ADDER_IN_from_mux[8][62] ,
         \ADDER_IN_from_mux[8][61] , \ADDER_IN_from_mux[8][60] ,
         \ADDER_IN_from_mux[8][59] , \ADDER_IN_from_mux[8][58] ,
         \ADDER_IN_from_mux[8][57] , \ADDER_IN_from_mux[8][56] ,
         \ADDER_IN_from_mux[8][55] , \ADDER_IN_from_mux[8][54] ,
         \ADDER_IN_from_mux[8][53] , \ADDER_IN_from_mux[8][52] ,
         \ADDER_IN_from_mux[8][51] , \ADDER_IN_from_mux[8][50] ,
         \ADDER_IN_from_mux[8][49] , \ADDER_IN_from_mux[8][48] ,
         \ADDER_IN_from_mux[8][47] , \ADDER_IN_from_mux[8][46] ,
         \ADDER_IN_from_mux[8][45] , \ADDER_IN_from_mux[8][44] ,
         \ADDER_IN_from_mux[8][43] , \ADDER_IN_from_mux[8][42] ,
         \ADDER_IN_from_mux[8][41] , \ADDER_IN_from_mux[8][40] ,
         \ADDER_IN_from_mux[8][39] , \ADDER_IN_from_mux[8][38] ,
         \ADDER_IN_from_mux[8][37] , \ADDER_IN_from_mux[8][36] ,
         \ADDER_IN_from_mux[8][35] , \ADDER_IN_from_mux[8][34] ,
         \ADDER_IN_from_mux[8][33] , \ADDER_IN_from_mux[8][32] ,
         \ADDER_IN_from_mux[8][31] , \ADDER_IN_from_mux[8][30] ,
         \ADDER_IN_from_mux[8][29] , \ADDER_IN_from_mux[8][28] ,
         \ADDER_IN_from_mux[8][27] , \ADDER_IN_from_mux[8][26] ,
         \ADDER_IN_from_mux[8][25] , \ADDER_IN_from_mux[8][24] ,
         \ADDER_IN_from_mux[8][23] , \ADDER_IN_from_mux[8][22] ,
         \ADDER_IN_from_mux[8][21] , \ADDER_IN_from_mux[8][20] ,
         \ADDER_IN_from_mux[8][19] , \ADDER_IN_from_mux[8][18] ,
         \ADDER_IN_from_mux[8][17] , \ADDER_IN_from_mux[8][16] ,
         \ADDER_IN_from_mux[8][15] , \ADDER_IN_from_mux[8][14] ,
         \ADDER_IN_from_mux[8][13] , \ADDER_IN_from_mux[8][12] ,
         \ADDER_IN_from_mux[8][11] , \ADDER_IN_from_mux[8][10] ,
         \ADDER_IN_from_mux[8][9] , \ADDER_IN_from_mux[8][8] ,
         \ADDER_IN_from_mux[8][7] , \ADDER_IN_from_mux[8][6] ,
         \ADDER_IN_from_mux[8][5] , \ADDER_IN_from_mux[8][4] ,
         \ADDER_IN_from_mux[8][3] , \ADDER_IN_from_mux[8][2] ,
         \ADDER_IN_from_mux[8][1] , \ADDER_IN_from_mux[8][0] ,
         \ADDER_IN_from_mux[7][63] , \ADDER_IN_from_mux[7][62] ,
         \ADDER_IN_from_mux[7][61] , \ADDER_IN_from_mux[7][60] ,
         \ADDER_IN_from_mux[7][59] , \ADDER_IN_from_mux[7][58] ,
         \ADDER_IN_from_mux[7][57] , \ADDER_IN_from_mux[7][56] ,
         \ADDER_IN_from_mux[7][55] , \ADDER_IN_from_mux[7][54] ,
         \ADDER_IN_from_mux[7][53] , \ADDER_IN_from_mux[7][52] ,
         \ADDER_IN_from_mux[7][51] , \ADDER_IN_from_mux[7][50] ,
         \ADDER_IN_from_mux[7][49] , \ADDER_IN_from_mux[7][48] ,
         \ADDER_IN_from_mux[7][47] , \ADDER_IN_from_mux[7][46] ,
         \ADDER_IN_from_mux[7][45] , \ADDER_IN_from_mux[7][44] ,
         \ADDER_IN_from_mux[7][43] , \ADDER_IN_from_mux[7][42] ,
         \ADDER_IN_from_mux[7][41] , \ADDER_IN_from_mux[7][40] ,
         \ADDER_IN_from_mux[7][39] , \ADDER_IN_from_mux[7][38] ,
         \ADDER_IN_from_mux[7][37] , \ADDER_IN_from_mux[7][36] ,
         \ADDER_IN_from_mux[7][35] , \ADDER_IN_from_mux[7][34] ,
         \ADDER_IN_from_mux[7][33] , \ADDER_IN_from_mux[7][32] ,
         \ADDER_IN_from_mux[7][31] , \ADDER_IN_from_mux[7][30] ,
         \ADDER_IN_from_mux[7][29] , \ADDER_IN_from_mux[7][28] ,
         \ADDER_IN_from_mux[7][27] , \ADDER_IN_from_mux[7][26] ,
         \ADDER_IN_from_mux[7][25] , \ADDER_IN_from_mux[7][24] ,
         \ADDER_IN_from_mux[7][23] , \ADDER_IN_from_mux[7][22] ,
         \ADDER_IN_from_mux[7][21] , \ADDER_IN_from_mux[7][20] ,
         \ADDER_IN_from_mux[7][19] , \ADDER_IN_from_mux[7][18] ,
         \ADDER_IN_from_mux[7][17] , \ADDER_IN_from_mux[7][16] ,
         \ADDER_IN_from_mux[7][15] , \ADDER_IN_from_mux[7][14] ,
         \ADDER_IN_from_mux[7][13] , \ADDER_IN_from_mux[7][12] ,
         \ADDER_IN_from_mux[7][11] , \ADDER_IN_from_mux[7][10] ,
         \ADDER_IN_from_mux[7][9] , \ADDER_IN_from_mux[7][8] ,
         \ADDER_IN_from_mux[7][7] , \ADDER_IN_from_mux[7][6] ,
         \ADDER_IN_from_mux[7][5] , \ADDER_IN_from_mux[7][4] ,
         \ADDER_IN_from_mux[7][3] , \ADDER_IN_from_mux[7][2] ,
         \ADDER_IN_from_mux[7][1] , \ADDER_IN_from_mux[7][0] ,
         \ADDER_IN_from_mux[6][63] , \ADDER_IN_from_mux[6][62] ,
         \ADDER_IN_from_mux[6][61] , \ADDER_IN_from_mux[6][60] ,
         \ADDER_IN_from_mux[6][59] , \ADDER_IN_from_mux[6][58] ,
         \ADDER_IN_from_mux[6][57] , \ADDER_IN_from_mux[6][56] ,
         \ADDER_IN_from_mux[6][55] , \ADDER_IN_from_mux[6][54] ,
         \ADDER_IN_from_mux[6][53] , \ADDER_IN_from_mux[6][52] ,
         \ADDER_IN_from_mux[6][51] , \ADDER_IN_from_mux[6][50] ,
         \ADDER_IN_from_mux[6][49] , \ADDER_IN_from_mux[6][48] ,
         \ADDER_IN_from_mux[6][47] , \ADDER_IN_from_mux[6][46] ,
         \ADDER_IN_from_mux[6][45] , \ADDER_IN_from_mux[6][44] ,
         \ADDER_IN_from_mux[6][43] , \ADDER_IN_from_mux[6][42] ,
         \ADDER_IN_from_mux[6][41] , \ADDER_IN_from_mux[6][40] ,
         \ADDER_IN_from_mux[6][39] , \ADDER_IN_from_mux[6][38] ,
         \ADDER_IN_from_mux[6][37] , \ADDER_IN_from_mux[6][36] ,
         \ADDER_IN_from_mux[6][35] , \ADDER_IN_from_mux[6][34] ,
         \ADDER_IN_from_mux[6][33] , \ADDER_IN_from_mux[6][32] ,
         \ADDER_IN_from_mux[6][31] , \ADDER_IN_from_mux[6][30] ,
         \ADDER_IN_from_mux[6][29] , \ADDER_IN_from_mux[6][28] ,
         \ADDER_IN_from_mux[6][27] , \ADDER_IN_from_mux[6][26] ,
         \ADDER_IN_from_mux[6][25] , \ADDER_IN_from_mux[6][24] ,
         \ADDER_IN_from_mux[6][23] , \ADDER_IN_from_mux[6][22] ,
         \ADDER_IN_from_mux[6][21] , \ADDER_IN_from_mux[6][20] ,
         \ADDER_IN_from_mux[6][19] , \ADDER_IN_from_mux[6][18] ,
         \ADDER_IN_from_mux[6][17] , \ADDER_IN_from_mux[6][16] ,
         \ADDER_IN_from_mux[6][15] , \ADDER_IN_from_mux[6][14] ,
         \ADDER_IN_from_mux[6][13] , \ADDER_IN_from_mux[6][12] ,
         \ADDER_IN_from_mux[6][11] , \ADDER_IN_from_mux[6][10] ,
         \ADDER_IN_from_mux[6][9] , \ADDER_IN_from_mux[6][8] ,
         \ADDER_IN_from_mux[6][7] , \ADDER_IN_from_mux[6][6] ,
         \ADDER_IN_from_mux[6][5] , \ADDER_IN_from_mux[6][4] ,
         \ADDER_IN_from_mux[6][3] , \ADDER_IN_from_mux[6][2] ,
         \ADDER_IN_from_mux[6][1] , \ADDER_IN_from_mux[6][0] ,
         \ADDER_IN_from_mux[5][63] , \ADDER_IN_from_mux[5][62] ,
         \ADDER_IN_from_mux[5][61] , \ADDER_IN_from_mux[5][60] ,
         \ADDER_IN_from_mux[5][59] , \ADDER_IN_from_mux[5][58] ,
         \ADDER_IN_from_mux[5][57] , \ADDER_IN_from_mux[5][56] ,
         \ADDER_IN_from_mux[5][55] , \ADDER_IN_from_mux[5][54] ,
         \ADDER_IN_from_mux[5][53] , \ADDER_IN_from_mux[5][52] ,
         \ADDER_IN_from_mux[5][51] , \ADDER_IN_from_mux[5][50] ,
         \ADDER_IN_from_mux[5][49] , \ADDER_IN_from_mux[5][48] ,
         \ADDER_IN_from_mux[5][47] , \ADDER_IN_from_mux[5][46] ,
         \ADDER_IN_from_mux[5][45] , \ADDER_IN_from_mux[5][44] ,
         \ADDER_IN_from_mux[5][43] , \ADDER_IN_from_mux[5][42] ,
         \ADDER_IN_from_mux[5][41] , \ADDER_IN_from_mux[5][40] ,
         \ADDER_IN_from_mux[5][39] , \ADDER_IN_from_mux[5][38] ,
         \ADDER_IN_from_mux[5][37] , \ADDER_IN_from_mux[5][36] ,
         \ADDER_IN_from_mux[5][35] , \ADDER_IN_from_mux[5][34] ,
         \ADDER_IN_from_mux[5][33] , \ADDER_IN_from_mux[5][32] ,
         \ADDER_IN_from_mux[5][31] , \ADDER_IN_from_mux[5][30] ,
         \ADDER_IN_from_mux[5][29] , \ADDER_IN_from_mux[5][28] ,
         \ADDER_IN_from_mux[5][27] , \ADDER_IN_from_mux[5][26] ,
         \ADDER_IN_from_mux[5][25] , \ADDER_IN_from_mux[5][24] ,
         \ADDER_IN_from_mux[5][23] , \ADDER_IN_from_mux[5][22] ,
         \ADDER_IN_from_mux[5][21] , \ADDER_IN_from_mux[5][20] ,
         \ADDER_IN_from_mux[5][19] , \ADDER_IN_from_mux[5][18] ,
         \ADDER_IN_from_mux[5][17] , \ADDER_IN_from_mux[5][16] ,
         \ADDER_IN_from_mux[5][15] , \ADDER_IN_from_mux[5][14] ,
         \ADDER_IN_from_mux[5][13] , \ADDER_IN_from_mux[5][12] ,
         \ADDER_IN_from_mux[5][11] , \ADDER_IN_from_mux[5][10] ,
         \ADDER_IN_from_mux[5][9] , \ADDER_IN_from_mux[5][8] ,
         \ADDER_IN_from_mux[5][7] , \ADDER_IN_from_mux[5][6] ,
         \ADDER_IN_from_mux[5][5] , \ADDER_IN_from_mux[5][4] ,
         \ADDER_IN_from_mux[5][3] , \ADDER_IN_from_mux[5][2] ,
         \ADDER_IN_from_mux[5][1] , \ADDER_IN_from_mux[5][0] ,
         \ADDER_IN_from_mux[4][63] , \ADDER_IN_from_mux[4][62] ,
         \ADDER_IN_from_mux[4][61] , \ADDER_IN_from_mux[4][60] ,
         \ADDER_IN_from_mux[4][59] , \ADDER_IN_from_mux[4][58] ,
         \ADDER_IN_from_mux[4][57] , \ADDER_IN_from_mux[4][56] ,
         \ADDER_IN_from_mux[4][55] , \ADDER_IN_from_mux[4][54] ,
         \ADDER_IN_from_mux[4][53] , \ADDER_IN_from_mux[4][52] ,
         \ADDER_IN_from_mux[4][51] , \ADDER_IN_from_mux[4][50] ,
         \ADDER_IN_from_mux[4][49] , \ADDER_IN_from_mux[4][48] ,
         \ADDER_IN_from_mux[4][47] , \ADDER_IN_from_mux[4][46] ,
         \ADDER_IN_from_mux[4][45] , \ADDER_IN_from_mux[4][44] ,
         \ADDER_IN_from_mux[4][43] , \ADDER_IN_from_mux[4][42] ,
         \ADDER_IN_from_mux[4][41] , \ADDER_IN_from_mux[4][40] ,
         \ADDER_IN_from_mux[4][39] , \ADDER_IN_from_mux[4][38] ,
         \ADDER_IN_from_mux[4][37] , \ADDER_IN_from_mux[4][36] ,
         \ADDER_IN_from_mux[4][35] , \ADDER_IN_from_mux[4][34] ,
         \ADDER_IN_from_mux[4][33] , \ADDER_IN_from_mux[4][32] ,
         \ADDER_IN_from_mux[4][31] , \ADDER_IN_from_mux[4][30] ,
         \ADDER_IN_from_mux[4][29] , \ADDER_IN_from_mux[4][28] ,
         \ADDER_IN_from_mux[4][27] , \ADDER_IN_from_mux[4][26] ,
         \ADDER_IN_from_mux[4][25] , \ADDER_IN_from_mux[4][24] ,
         \ADDER_IN_from_mux[4][23] , \ADDER_IN_from_mux[4][22] ,
         \ADDER_IN_from_mux[4][21] , \ADDER_IN_from_mux[4][20] ,
         \ADDER_IN_from_mux[4][19] , \ADDER_IN_from_mux[4][18] ,
         \ADDER_IN_from_mux[4][17] , \ADDER_IN_from_mux[4][16] ,
         \ADDER_IN_from_mux[4][15] , \ADDER_IN_from_mux[4][14] ,
         \ADDER_IN_from_mux[4][13] , \ADDER_IN_from_mux[4][12] ,
         \ADDER_IN_from_mux[4][11] , \ADDER_IN_from_mux[4][10] ,
         \ADDER_IN_from_mux[4][9] , \ADDER_IN_from_mux[4][8] ,
         \ADDER_IN_from_mux[4][7] , \ADDER_IN_from_mux[4][6] ,
         \ADDER_IN_from_mux[4][5] , \ADDER_IN_from_mux[4][4] ,
         \ADDER_IN_from_mux[4][3] , \ADDER_IN_from_mux[4][2] ,
         \ADDER_IN_from_mux[4][1] , \ADDER_IN_from_mux[4][0] ,
         \ADDER_IN_from_mux[3][63] , \ADDER_IN_from_mux[3][62] ,
         \ADDER_IN_from_mux[3][61] , \ADDER_IN_from_mux[3][60] ,
         \ADDER_IN_from_mux[3][59] , \ADDER_IN_from_mux[3][58] ,
         \ADDER_IN_from_mux[3][57] , \ADDER_IN_from_mux[3][56] ,
         \ADDER_IN_from_mux[3][55] , \ADDER_IN_from_mux[3][54] ,
         \ADDER_IN_from_mux[3][53] , \ADDER_IN_from_mux[3][52] ,
         \ADDER_IN_from_mux[3][51] , \ADDER_IN_from_mux[3][50] ,
         \ADDER_IN_from_mux[3][49] , \ADDER_IN_from_mux[3][48] ,
         \ADDER_IN_from_mux[3][47] , \ADDER_IN_from_mux[3][46] ,
         \ADDER_IN_from_mux[3][45] , \ADDER_IN_from_mux[3][44] ,
         \ADDER_IN_from_mux[3][43] , \ADDER_IN_from_mux[3][42] ,
         \ADDER_IN_from_mux[3][41] , \ADDER_IN_from_mux[3][40] ,
         \ADDER_IN_from_mux[3][39] , \ADDER_IN_from_mux[3][38] ,
         \ADDER_IN_from_mux[3][37] , \ADDER_IN_from_mux[3][36] ,
         \ADDER_IN_from_mux[3][35] , \ADDER_IN_from_mux[3][34] ,
         \ADDER_IN_from_mux[3][33] , \ADDER_IN_from_mux[3][32] ,
         \ADDER_IN_from_mux[3][31] , \ADDER_IN_from_mux[3][30] ,
         \ADDER_IN_from_mux[3][29] , \ADDER_IN_from_mux[3][28] ,
         \ADDER_IN_from_mux[3][27] , \ADDER_IN_from_mux[3][26] ,
         \ADDER_IN_from_mux[3][25] , \ADDER_IN_from_mux[3][24] ,
         \ADDER_IN_from_mux[3][23] , \ADDER_IN_from_mux[3][22] ,
         \ADDER_IN_from_mux[3][21] , \ADDER_IN_from_mux[3][20] ,
         \ADDER_IN_from_mux[3][19] , \ADDER_IN_from_mux[3][18] ,
         \ADDER_IN_from_mux[3][17] , \ADDER_IN_from_mux[3][16] ,
         \ADDER_IN_from_mux[3][15] , \ADDER_IN_from_mux[3][14] ,
         \ADDER_IN_from_mux[3][13] , \ADDER_IN_from_mux[3][12] ,
         \ADDER_IN_from_mux[3][11] , \ADDER_IN_from_mux[3][10] ,
         \ADDER_IN_from_mux[3][9] , \ADDER_IN_from_mux[3][8] ,
         \ADDER_IN_from_mux[3][7] , \ADDER_IN_from_mux[3][6] ,
         \ADDER_IN_from_mux[3][5] , \ADDER_IN_from_mux[3][4] ,
         \ADDER_IN_from_mux[3][3] , \ADDER_IN_from_mux[3][2] ,
         \ADDER_IN_from_mux[3][1] , \ADDER_IN_from_mux[3][0] ,
         \ADDER_IN_from_mux[2][63] , \ADDER_IN_from_mux[2][62] ,
         \ADDER_IN_from_mux[2][61] , \ADDER_IN_from_mux[2][60] ,
         \ADDER_IN_from_mux[2][59] , \ADDER_IN_from_mux[2][58] ,
         \ADDER_IN_from_mux[2][57] , \ADDER_IN_from_mux[2][56] ,
         \ADDER_IN_from_mux[2][55] , \ADDER_IN_from_mux[2][54] ,
         \ADDER_IN_from_mux[2][53] , \ADDER_IN_from_mux[2][52] ,
         \ADDER_IN_from_mux[2][51] , \ADDER_IN_from_mux[2][50] ,
         \ADDER_IN_from_mux[2][49] , \ADDER_IN_from_mux[2][48] ,
         \ADDER_IN_from_mux[2][47] , \ADDER_IN_from_mux[2][46] ,
         \ADDER_IN_from_mux[2][45] , \ADDER_IN_from_mux[2][44] ,
         \ADDER_IN_from_mux[2][43] , \ADDER_IN_from_mux[2][42] ,
         \ADDER_IN_from_mux[2][41] , \ADDER_IN_from_mux[2][40] ,
         \ADDER_IN_from_mux[2][39] , \ADDER_IN_from_mux[2][38] ,
         \ADDER_IN_from_mux[2][37] , \ADDER_IN_from_mux[2][36] ,
         \ADDER_IN_from_mux[2][35] , \ADDER_IN_from_mux[2][34] ,
         \ADDER_IN_from_mux[2][33] , \ADDER_IN_from_mux[2][32] ,
         \ADDER_IN_from_mux[2][31] , \ADDER_IN_from_mux[2][30] ,
         \ADDER_IN_from_mux[2][29] , \ADDER_IN_from_mux[2][28] ,
         \ADDER_IN_from_mux[2][27] , \ADDER_IN_from_mux[2][26] ,
         \ADDER_IN_from_mux[2][25] , \ADDER_IN_from_mux[2][24] ,
         \ADDER_IN_from_mux[2][23] , \ADDER_IN_from_mux[2][22] ,
         \ADDER_IN_from_mux[2][21] , \ADDER_IN_from_mux[2][20] ,
         \ADDER_IN_from_mux[2][19] , \ADDER_IN_from_mux[2][18] ,
         \ADDER_IN_from_mux[2][17] , \ADDER_IN_from_mux[2][16] ,
         \ADDER_IN_from_mux[2][15] , \ADDER_IN_from_mux[2][14] ,
         \ADDER_IN_from_mux[2][13] , \ADDER_IN_from_mux[2][12] ,
         \ADDER_IN_from_mux[2][11] , \ADDER_IN_from_mux[2][10] ,
         \ADDER_IN_from_mux[2][9] , \ADDER_IN_from_mux[2][8] ,
         \ADDER_IN_from_mux[2][7] , \ADDER_IN_from_mux[2][6] ,
         \ADDER_IN_from_mux[2][5] , \ADDER_IN_from_mux[2][4] ,
         \ADDER_IN_from_mux[2][3] , \ADDER_IN_from_mux[2][2] ,
         \ADDER_IN_from_mux[2][1] , \ADDER_IN_from_mux[2][0] ,
         \ADDER_IN_from_mux[1][63] , \ADDER_IN_from_mux[1][62] ,
         \ADDER_IN_from_mux[1][61] , \ADDER_IN_from_mux[1][60] ,
         \ADDER_IN_from_mux[1][59] , \ADDER_IN_from_mux[1][58] ,
         \ADDER_IN_from_mux[1][57] , \ADDER_IN_from_mux[1][56] ,
         \ADDER_IN_from_mux[1][55] , \ADDER_IN_from_mux[1][54] ,
         \ADDER_IN_from_mux[1][53] , \ADDER_IN_from_mux[1][52] ,
         \ADDER_IN_from_mux[1][51] , \ADDER_IN_from_mux[1][50] ,
         \ADDER_IN_from_mux[1][49] , \ADDER_IN_from_mux[1][48] ,
         \ADDER_IN_from_mux[1][47] , \ADDER_IN_from_mux[1][46] ,
         \ADDER_IN_from_mux[1][45] , \ADDER_IN_from_mux[1][44] ,
         \ADDER_IN_from_mux[1][43] , \ADDER_IN_from_mux[1][42] ,
         \ADDER_IN_from_mux[1][41] , \ADDER_IN_from_mux[1][40] ,
         \ADDER_IN_from_mux[1][39] , \ADDER_IN_from_mux[1][38] ,
         \ADDER_IN_from_mux[1][37] , \ADDER_IN_from_mux[1][36] ,
         \ADDER_IN_from_mux[1][35] , \ADDER_IN_from_mux[1][34] ,
         \ADDER_IN_from_mux[1][33] , \ADDER_IN_from_mux[1][32] ,
         \ADDER_IN_from_mux[1][31] , \ADDER_IN_from_mux[1][30] ,
         \ADDER_IN_from_mux[1][29] , \ADDER_IN_from_mux[1][28] ,
         \ADDER_IN_from_mux[1][27] , \ADDER_IN_from_mux[1][26] ,
         \ADDER_IN_from_mux[1][25] , \ADDER_IN_from_mux[1][24] ,
         \ADDER_IN_from_mux[1][23] , \ADDER_IN_from_mux[1][22] ,
         \ADDER_IN_from_mux[1][21] , \ADDER_IN_from_mux[1][20] ,
         \ADDER_IN_from_mux[1][19] , \ADDER_IN_from_mux[1][18] ,
         \ADDER_IN_from_mux[1][17] , \ADDER_IN_from_mux[1][16] ,
         \ADDER_IN_from_mux[1][15] , \ADDER_IN_from_mux[1][14] ,
         \ADDER_IN_from_mux[1][13] , \ADDER_IN_from_mux[1][12] ,
         \ADDER_IN_from_mux[1][11] , \ADDER_IN_from_mux[1][10] ,
         \ADDER_IN_from_mux[1][9] , \ADDER_IN_from_mux[1][8] ,
         \ADDER_IN_from_mux[1][7] , \ADDER_IN_from_mux[1][6] ,
         \ADDER_IN_from_mux[1][5] , \ADDER_IN_from_mux[1][4] ,
         \ADDER_IN_from_mux[1][3] , \ADDER_IN_from_mux[1][2] ,
         \ADDER_IN_from_mux[1][1] , \ADDER_IN_from_mux[1][0] ,
         \ADDER_IN_from_mux[0][63] , \ADDER_IN_from_mux[0][62] ,
         \ADDER_IN_from_mux[0][61] , \ADDER_IN_from_mux[0][60] ,
         \ADDER_IN_from_mux[0][59] , \ADDER_IN_from_mux[0][58] ,
         \ADDER_IN_from_mux[0][57] , \ADDER_IN_from_mux[0][56] ,
         \ADDER_IN_from_mux[0][55] , \ADDER_IN_from_mux[0][54] ,
         \ADDER_IN_from_mux[0][53] , \ADDER_IN_from_mux[0][52] ,
         \ADDER_IN_from_mux[0][51] , \ADDER_IN_from_mux[0][50] ,
         \ADDER_IN_from_mux[0][49] , \ADDER_IN_from_mux[0][48] ,
         \ADDER_IN_from_mux[0][47] , \ADDER_IN_from_mux[0][46] ,
         \ADDER_IN_from_mux[0][45] , \ADDER_IN_from_mux[0][44] ,
         \ADDER_IN_from_mux[0][43] , \ADDER_IN_from_mux[0][42] ,
         \ADDER_IN_from_mux[0][41] , \ADDER_IN_from_mux[0][40] ,
         \ADDER_IN_from_mux[0][39] , \ADDER_IN_from_mux[0][38] ,
         \ADDER_IN_from_mux[0][37] , \ADDER_IN_from_mux[0][36] ,
         \ADDER_IN_from_mux[0][35] , \ADDER_IN_from_mux[0][34] ,
         \ADDER_IN_from_mux[0][33] , \ADDER_IN_from_mux[0][32] ,
         \ADDER_IN_from_mux[0][31] , \ADDER_IN_from_mux[0][30] ,
         \ADDER_IN_from_mux[0][29] , \ADDER_IN_from_mux[0][28] ,
         \ADDER_IN_from_mux[0][27] , \ADDER_IN_from_mux[0][26] ,
         \ADDER_IN_from_mux[0][25] , \ADDER_IN_from_mux[0][24] ,
         \ADDER_IN_from_mux[0][23] , \ADDER_IN_from_mux[0][22] ,
         \ADDER_IN_from_mux[0][21] , \ADDER_IN_from_mux[0][20] ,
         \ADDER_IN_from_mux[0][19] , \ADDER_IN_from_mux[0][18] ,
         \ADDER_IN_from_mux[0][17] , \ADDER_IN_from_mux[0][16] ,
         \ADDER_IN_from_mux[0][15] , \ADDER_IN_from_mux[0][14] ,
         \ADDER_IN_from_mux[0][13] , \ADDER_IN_from_mux[0][12] ,
         \ADDER_IN_from_mux[0][11] , \ADDER_IN_from_mux[0][10] ,
         \ADDER_IN_from_mux[0][9] , \ADDER_IN_from_mux[0][8] ,
         \ADDER_IN_from_mux[0][7] , \ADDER_IN_from_mux[0][6] ,
         \ADDER_IN_from_mux[0][5] , \ADDER_IN_from_mux[0][4] ,
         \ADDER_IN_from_mux[0][3] , \ADDER_IN_from_mux[0][2] ,
         \ADDER_IN_from_mux[0][1] , \ADDER_IN_from_mux[0][0] ,
         \ADDER_IN_from_sum[14][63] , \ADDER_IN_from_sum[14][62] ,
         \ADDER_IN_from_sum[14][61] , \ADDER_IN_from_sum[14][60] ,
         \ADDER_IN_from_sum[14][59] , \ADDER_IN_from_sum[14][58] ,
         \ADDER_IN_from_sum[14][57] , \ADDER_IN_from_sum[14][56] ,
         \ADDER_IN_from_sum[14][55] , \ADDER_IN_from_sum[14][54] ,
         \ADDER_IN_from_sum[14][53] , \ADDER_IN_from_sum[14][52] ,
         \ADDER_IN_from_sum[14][51] , \ADDER_IN_from_sum[14][50] ,
         \ADDER_IN_from_sum[14][49] , \ADDER_IN_from_sum[14][48] ,
         \ADDER_IN_from_sum[14][47] , \ADDER_IN_from_sum[14][46] ,
         \ADDER_IN_from_sum[14][45] , \ADDER_IN_from_sum[14][44] ,
         \ADDER_IN_from_sum[14][43] , \ADDER_IN_from_sum[14][42] ,
         \ADDER_IN_from_sum[14][41] , \ADDER_IN_from_sum[14][40] ,
         \ADDER_IN_from_sum[14][39] , \ADDER_IN_from_sum[14][38] ,
         \ADDER_IN_from_sum[14][37] , \ADDER_IN_from_sum[14][36] ,
         \ADDER_IN_from_sum[14][35] , \ADDER_IN_from_sum[14][34] ,
         \ADDER_IN_from_sum[14][33] , \ADDER_IN_from_sum[14][32] ,
         \ADDER_IN_from_sum[14][31] , \ADDER_IN_from_sum[14][30] ,
         \ADDER_IN_from_sum[14][29] , \ADDER_IN_from_sum[14][28] ,
         \ADDER_IN_from_sum[14][27] , \ADDER_IN_from_sum[14][26] ,
         \ADDER_IN_from_sum[14][25] , \ADDER_IN_from_sum[14][24] ,
         \ADDER_IN_from_sum[14][23] , \ADDER_IN_from_sum[14][22] ,
         \ADDER_IN_from_sum[14][21] , \ADDER_IN_from_sum[14][20] ,
         \ADDER_IN_from_sum[14][19] , \ADDER_IN_from_sum[14][18] ,
         \ADDER_IN_from_sum[14][17] , \ADDER_IN_from_sum[14][16] ,
         \ADDER_IN_from_sum[14][15] , \ADDER_IN_from_sum[14][14] ,
         \ADDER_IN_from_sum[14][13] , \ADDER_IN_from_sum[14][12] ,
         \ADDER_IN_from_sum[14][11] , \ADDER_IN_from_sum[14][10] ,
         \ADDER_IN_from_sum[14][9] , \ADDER_IN_from_sum[14][8] ,
         \ADDER_IN_from_sum[14][7] , \ADDER_IN_from_sum[14][6] ,
         \ADDER_IN_from_sum[14][5] , \ADDER_IN_from_sum[14][4] ,
         \ADDER_IN_from_sum[14][3] , \ADDER_IN_from_sum[14][2] ,
         \ADDER_IN_from_sum[14][1] , \ADDER_IN_from_sum[14][0] ,
         \ADDER_IN_from_sum[13][63] , \ADDER_IN_from_sum[13][62] ,
         \ADDER_IN_from_sum[13][61] , \ADDER_IN_from_sum[13][60] ,
         \ADDER_IN_from_sum[13][59] , \ADDER_IN_from_sum[13][58] ,
         \ADDER_IN_from_sum[13][57] , \ADDER_IN_from_sum[13][56] ,
         \ADDER_IN_from_sum[13][55] , \ADDER_IN_from_sum[13][54] ,
         \ADDER_IN_from_sum[13][53] , \ADDER_IN_from_sum[13][52] ,
         \ADDER_IN_from_sum[13][51] , \ADDER_IN_from_sum[13][50] ,
         \ADDER_IN_from_sum[13][49] , \ADDER_IN_from_sum[13][48] ,
         \ADDER_IN_from_sum[13][47] , \ADDER_IN_from_sum[13][46] ,
         \ADDER_IN_from_sum[13][45] , \ADDER_IN_from_sum[13][44] ,
         \ADDER_IN_from_sum[13][43] , \ADDER_IN_from_sum[13][42] ,
         \ADDER_IN_from_sum[13][41] , \ADDER_IN_from_sum[13][40] ,
         \ADDER_IN_from_sum[13][39] , \ADDER_IN_from_sum[13][38] ,
         \ADDER_IN_from_sum[13][37] , \ADDER_IN_from_sum[13][36] ,
         \ADDER_IN_from_sum[13][35] , \ADDER_IN_from_sum[13][34] ,
         \ADDER_IN_from_sum[13][33] , \ADDER_IN_from_sum[13][32] ,
         \ADDER_IN_from_sum[13][31] , \ADDER_IN_from_sum[13][30] ,
         \ADDER_IN_from_sum[13][29] , \ADDER_IN_from_sum[13][28] ,
         \ADDER_IN_from_sum[13][27] , \ADDER_IN_from_sum[13][26] ,
         \ADDER_IN_from_sum[13][25] , \ADDER_IN_from_sum[13][24] ,
         \ADDER_IN_from_sum[13][23] , \ADDER_IN_from_sum[13][22] ,
         \ADDER_IN_from_sum[13][21] , \ADDER_IN_from_sum[13][20] ,
         \ADDER_IN_from_sum[13][19] , \ADDER_IN_from_sum[13][18] ,
         \ADDER_IN_from_sum[13][17] , \ADDER_IN_from_sum[13][16] ,
         \ADDER_IN_from_sum[13][15] , \ADDER_IN_from_sum[13][14] ,
         \ADDER_IN_from_sum[13][13] , \ADDER_IN_from_sum[13][12] ,
         \ADDER_IN_from_sum[13][11] , \ADDER_IN_from_sum[13][10] ,
         \ADDER_IN_from_sum[13][9] , \ADDER_IN_from_sum[13][8] ,
         \ADDER_IN_from_sum[13][7] , \ADDER_IN_from_sum[13][6] ,
         \ADDER_IN_from_sum[13][5] , \ADDER_IN_from_sum[13][4] ,
         \ADDER_IN_from_sum[13][3] , \ADDER_IN_from_sum[13][2] ,
         \ADDER_IN_from_sum[13][1] , \ADDER_IN_from_sum[13][0] ,
         \ADDER_IN_from_sum[12][63] , \ADDER_IN_from_sum[12][62] ,
         \ADDER_IN_from_sum[12][61] , \ADDER_IN_from_sum[12][60] ,
         \ADDER_IN_from_sum[12][59] , \ADDER_IN_from_sum[12][58] ,
         \ADDER_IN_from_sum[12][57] , \ADDER_IN_from_sum[12][56] ,
         \ADDER_IN_from_sum[12][55] , \ADDER_IN_from_sum[12][54] ,
         \ADDER_IN_from_sum[12][53] , \ADDER_IN_from_sum[12][52] ,
         \ADDER_IN_from_sum[12][51] , \ADDER_IN_from_sum[12][50] ,
         \ADDER_IN_from_sum[12][49] , \ADDER_IN_from_sum[12][48] ,
         \ADDER_IN_from_sum[12][47] , \ADDER_IN_from_sum[12][46] ,
         \ADDER_IN_from_sum[12][45] , \ADDER_IN_from_sum[12][44] ,
         \ADDER_IN_from_sum[12][43] , \ADDER_IN_from_sum[12][42] ,
         \ADDER_IN_from_sum[12][41] , \ADDER_IN_from_sum[12][40] ,
         \ADDER_IN_from_sum[12][39] , \ADDER_IN_from_sum[12][38] ,
         \ADDER_IN_from_sum[12][37] , \ADDER_IN_from_sum[12][36] ,
         \ADDER_IN_from_sum[12][35] , \ADDER_IN_from_sum[12][34] ,
         \ADDER_IN_from_sum[12][33] , \ADDER_IN_from_sum[12][32] ,
         \ADDER_IN_from_sum[12][31] , \ADDER_IN_from_sum[12][30] ,
         \ADDER_IN_from_sum[12][29] , \ADDER_IN_from_sum[12][28] ,
         \ADDER_IN_from_sum[12][27] , \ADDER_IN_from_sum[12][26] ,
         \ADDER_IN_from_sum[12][25] , \ADDER_IN_from_sum[12][24] ,
         \ADDER_IN_from_sum[12][23] , \ADDER_IN_from_sum[12][22] ,
         \ADDER_IN_from_sum[12][21] , \ADDER_IN_from_sum[12][20] ,
         \ADDER_IN_from_sum[12][19] , \ADDER_IN_from_sum[12][18] ,
         \ADDER_IN_from_sum[12][17] , \ADDER_IN_from_sum[12][16] ,
         \ADDER_IN_from_sum[12][15] , \ADDER_IN_from_sum[12][14] ,
         \ADDER_IN_from_sum[12][13] , \ADDER_IN_from_sum[12][12] ,
         \ADDER_IN_from_sum[12][11] , \ADDER_IN_from_sum[12][10] ,
         \ADDER_IN_from_sum[12][9] , \ADDER_IN_from_sum[12][8] ,
         \ADDER_IN_from_sum[12][7] , \ADDER_IN_from_sum[12][6] ,
         \ADDER_IN_from_sum[12][5] , \ADDER_IN_from_sum[12][4] ,
         \ADDER_IN_from_sum[12][3] , \ADDER_IN_from_sum[12][2] ,
         \ADDER_IN_from_sum[12][1] , \ADDER_IN_from_sum[12][0] ,
         \ADDER_IN_from_sum[11][63] , \ADDER_IN_from_sum[11][62] ,
         \ADDER_IN_from_sum[11][61] , \ADDER_IN_from_sum[11][60] ,
         \ADDER_IN_from_sum[11][59] , \ADDER_IN_from_sum[11][58] ,
         \ADDER_IN_from_sum[11][57] , \ADDER_IN_from_sum[11][56] ,
         \ADDER_IN_from_sum[11][55] , \ADDER_IN_from_sum[11][54] ,
         \ADDER_IN_from_sum[11][53] , \ADDER_IN_from_sum[11][52] ,
         \ADDER_IN_from_sum[11][51] , \ADDER_IN_from_sum[11][50] ,
         \ADDER_IN_from_sum[11][49] , \ADDER_IN_from_sum[11][48] ,
         \ADDER_IN_from_sum[11][47] , \ADDER_IN_from_sum[11][46] ,
         \ADDER_IN_from_sum[11][45] , \ADDER_IN_from_sum[11][44] ,
         \ADDER_IN_from_sum[11][43] , \ADDER_IN_from_sum[11][42] ,
         \ADDER_IN_from_sum[11][41] , \ADDER_IN_from_sum[11][40] ,
         \ADDER_IN_from_sum[11][39] , \ADDER_IN_from_sum[11][38] ,
         \ADDER_IN_from_sum[11][37] , \ADDER_IN_from_sum[11][36] ,
         \ADDER_IN_from_sum[11][35] , \ADDER_IN_from_sum[11][34] ,
         \ADDER_IN_from_sum[11][33] , \ADDER_IN_from_sum[11][32] ,
         \ADDER_IN_from_sum[11][31] , \ADDER_IN_from_sum[11][30] ,
         \ADDER_IN_from_sum[11][29] , \ADDER_IN_from_sum[11][28] ,
         \ADDER_IN_from_sum[11][27] , \ADDER_IN_from_sum[11][26] ,
         \ADDER_IN_from_sum[11][25] , \ADDER_IN_from_sum[11][24] ,
         \ADDER_IN_from_sum[11][23] , \ADDER_IN_from_sum[11][22] ,
         \ADDER_IN_from_sum[11][21] , \ADDER_IN_from_sum[11][20] ,
         \ADDER_IN_from_sum[11][19] , \ADDER_IN_from_sum[11][18] ,
         \ADDER_IN_from_sum[11][17] , \ADDER_IN_from_sum[11][16] ,
         \ADDER_IN_from_sum[11][15] , \ADDER_IN_from_sum[11][14] ,
         \ADDER_IN_from_sum[11][13] , \ADDER_IN_from_sum[11][12] ,
         \ADDER_IN_from_sum[11][11] , \ADDER_IN_from_sum[11][10] ,
         \ADDER_IN_from_sum[11][9] , \ADDER_IN_from_sum[11][8] ,
         \ADDER_IN_from_sum[11][7] , \ADDER_IN_from_sum[11][6] ,
         \ADDER_IN_from_sum[11][5] , \ADDER_IN_from_sum[11][4] ,
         \ADDER_IN_from_sum[11][3] , \ADDER_IN_from_sum[11][2] ,
         \ADDER_IN_from_sum[11][1] , \ADDER_IN_from_sum[11][0] ,
         \ADDER_IN_from_sum[10][63] , \ADDER_IN_from_sum[10][62] ,
         \ADDER_IN_from_sum[10][61] , \ADDER_IN_from_sum[10][60] ,
         \ADDER_IN_from_sum[10][59] , \ADDER_IN_from_sum[10][58] ,
         \ADDER_IN_from_sum[10][57] , \ADDER_IN_from_sum[10][56] ,
         \ADDER_IN_from_sum[10][55] , \ADDER_IN_from_sum[10][54] ,
         \ADDER_IN_from_sum[10][53] , \ADDER_IN_from_sum[10][52] ,
         \ADDER_IN_from_sum[10][51] , \ADDER_IN_from_sum[10][50] ,
         \ADDER_IN_from_sum[10][49] , \ADDER_IN_from_sum[10][48] ,
         \ADDER_IN_from_sum[10][47] , \ADDER_IN_from_sum[10][46] ,
         \ADDER_IN_from_sum[10][45] , \ADDER_IN_from_sum[10][44] ,
         \ADDER_IN_from_sum[10][43] , \ADDER_IN_from_sum[10][42] ,
         \ADDER_IN_from_sum[10][41] , \ADDER_IN_from_sum[10][40] ,
         \ADDER_IN_from_sum[10][39] , \ADDER_IN_from_sum[10][38] ,
         \ADDER_IN_from_sum[10][37] , \ADDER_IN_from_sum[10][36] ,
         \ADDER_IN_from_sum[10][35] , \ADDER_IN_from_sum[10][34] ,
         \ADDER_IN_from_sum[10][33] , \ADDER_IN_from_sum[10][32] ,
         \ADDER_IN_from_sum[10][31] , \ADDER_IN_from_sum[10][30] ,
         \ADDER_IN_from_sum[10][29] , \ADDER_IN_from_sum[10][28] ,
         \ADDER_IN_from_sum[10][27] , \ADDER_IN_from_sum[10][26] ,
         \ADDER_IN_from_sum[10][25] , \ADDER_IN_from_sum[10][24] ,
         \ADDER_IN_from_sum[10][23] , \ADDER_IN_from_sum[10][22] ,
         \ADDER_IN_from_sum[10][21] , \ADDER_IN_from_sum[10][20] ,
         \ADDER_IN_from_sum[10][19] , \ADDER_IN_from_sum[10][18] ,
         \ADDER_IN_from_sum[10][17] , \ADDER_IN_from_sum[10][16] ,
         \ADDER_IN_from_sum[10][15] , \ADDER_IN_from_sum[10][14] ,
         \ADDER_IN_from_sum[10][13] , \ADDER_IN_from_sum[10][12] ,
         \ADDER_IN_from_sum[10][11] , \ADDER_IN_from_sum[10][10] ,
         \ADDER_IN_from_sum[10][9] , \ADDER_IN_from_sum[10][8] ,
         \ADDER_IN_from_sum[10][7] , \ADDER_IN_from_sum[10][6] ,
         \ADDER_IN_from_sum[10][5] , \ADDER_IN_from_sum[10][4] ,
         \ADDER_IN_from_sum[10][3] , \ADDER_IN_from_sum[10][2] ,
         \ADDER_IN_from_sum[10][1] , \ADDER_IN_from_sum[10][0] ,
         \ADDER_IN_from_sum[9][63] , \ADDER_IN_from_sum[9][62] ,
         \ADDER_IN_from_sum[9][61] , \ADDER_IN_from_sum[9][60] ,
         \ADDER_IN_from_sum[9][59] , \ADDER_IN_from_sum[9][58] ,
         \ADDER_IN_from_sum[9][57] , \ADDER_IN_from_sum[9][56] ,
         \ADDER_IN_from_sum[9][55] , \ADDER_IN_from_sum[9][54] ,
         \ADDER_IN_from_sum[9][53] , \ADDER_IN_from_sum[9][52] ,
         \ADDER_IN_from_sum[9][51] , \ADDER_IN_from_sum[9][50] ,
         \ADDER_IN_from_sum[9][49] , \ADDER_IN_from_sum[9][48] ,
         \ADDER_IN_from_sum[9][47] , \ADDER_IN_from_sum[9][46] ,
         \ADDER_IN_from_sum[9][45] , \ADDER_IN_from_sum[9][44] ,
         \ADDER_IN_from_sum[9][43] , \ADDER_IN_from_sum[9][42] ,
         \ADDER_IN_from_sum[9][41] , \ADDER_IN_from_sum[9][40] ,
         \ADDER_IN_from_sum[9][39] , \ADDER_IN_from_sum[9][38] ,
         \ADDER_IN_from_sum[9][37] , \ADDER_IN_from_sum[9][36] ,
         \ADDER_IN_from_sum[9][35] , \ADDER_IN_from_sum[9][34] ,
         \ADDER_IN_from_sum[9][33] , \ADDER_IN_from_sum[9][32] ,
         \ADDER_IN_from_sum[9][31] , \ADDER_IN_from_sum[9][30] ,
         \ADDER_IN_from_sum[9][29] , \ADDER_IN_from_sum[9][28] ,
         \ADDER_IN_from_sum[9][27] , \ADDER_IN_from_sum[9][26] ,
         \ADDER_IN_from_sum[9][25] , \ADDER_IN_from_sum[9][24] ,
         \ADDER_IN_from_sum[9][23] , \ADDER_IN_from_sum[9][22] ,
         \ADDER_IN_from_sum[9][21] , \ADDER_IN_from_sum[9][20] ,
         \ADDER_IN_from_sum[9][19] , \ADDER_IN_from_sum[9][18] ,
         \ADDER_IN_from_sum[9][17] , \ADDER_IN_from_sum[9][16] ,
         \ADDER_IN_from_sum[9][15] , \ADDER_IN_from_sum[9][14] ,
         \ADDER_IN_from_sum[9][13] , \ADDER_IN_from_sum[9][12] ,
         \ADDER_IN_from_sum[9][11] , \ADDER_IN_from_sum[9][10] ,
         \ADDER_IN_from_sum[9][9] , \ADDER_IN_from_sum[9][8] ,
         \ADDER_IN_from_sum[9][7] , \ADDER_IN_from_sum[9][6] ,
         \ADDER_IN_from_sum[9][5] , \ADDER_IN_from_sum[9][4] ,
         \ADDER_IN_from_sum[9][3] , \ADDER_IN_from_sum[9][2] ,
         \ADDER_IN_from_sum[9][1] , \ADDER_IN_from_sum[9][0] ,
         \ADDER_IN_from_sum[8][63] , \ADDER_IN_from_sum[8][62] ,
         \ADDER_IN_from_sum[8][61] , \ADDER_IN_from_sum[8][60] ,
         \ADDER_IN_from_sum[8][59] , \ADDER_IN_from_sum[8][58] ,
         \ADDER_IN_from_sum[8][57] , \ADDER_IN_from_sum[8][56] ,
         \ADDER_IN_from_sum[8][55] , \ADDER_IN_from_sum[8][54] ,
         \ADDER_IN_from_sum[8][53] , \ADDER_IN_from_sum[8][52] ,
         \ADDER_IN_from_sum[8][51] , \ADDER_IN_from_sum[8][50] ,
         \ADDER_IN_from_sum[8][49] , \ADDER_IN_from_sum[8][48] ,
         \ADDER_IN_from_sum[8][47] , \ADDER_IN_from_sum[8][46] ,
         \ADDER_IN_from_sum[8][45] , \ADDER_IN_from_sum[8][44] ,
         \ADDER_IN_from_sum[8][43] , \ADDER_IN_from_sum[8][42] ,
         \ADDER_IN_from_sum[8][41] , \ADDER_IN_from_sum[8][40] ,
         \ADDER_IN_from_sum[8][39] , \ADDER_IN_from_sum[8][38] ,
         \ADDER_IN_from_sum[8][37] , \ADDER_IN_from_sum[8][36] ,
         \ADDER_IN_from_sum[8][35] , \ADDER_IN_from_sum[8][34] ,
         \ADDER_IN_from_sum[8][33] , \ADDER_IN_from_sum[8][32] ,
         \ADDER_IN_from_sum[8][31] , \ADDER_IN_from_sum[8][30] ,
         \ADDER_IN_from_sum[8][29] , \ADDER_IN_from_sum[8][28] ,
         \ADDER_IN_from_sum[8][27] , \ADDER_IN_from_sum[8][26] ,
         \ADDER_IN_from_sum[8][25] , \ADDER_IN_from_sum[8][24] ,
         \ADDER_IN_from_sum[8][23] , \ADDER_IN_from_sum[8][22] ,
         \ADDER_IN_from_sum[8][21] , \ADDER_IN_from_sum[8][20] ,
         \ADDER_IN_from_sum[8][19] , \ADDER_IN_from_sum[8][18] ,
         \ADDER_IN_from_sum[8][17] , \ADDER_IN_from_sum[8][16] ,
         \ADDER_IN_from_sum[8][15] , \ADDER_IN_from_sum[8][14] ,
         \ADDER_IN_from_sum[8][13] , \ADDER_IN_from_sum[8][12] ,
         \ADDER_IN_from_sum[8][11] , \ADDER_IN_from_sum[8][10] ,
         \ADDER_IN_from_sum[8][9] , \ADDER_IN_from_sum[8][8] ,
         \ADDER_IN_from_sum[8][7] , \ADDER_IN_from_sum[8][6] ,
         \ADDER_IN_from_sum[8][5] , \ADDER_IN_from_sum[8][4] ,
         \ADDER_IN_from_sum[8][3] , \ADDER_IN_from_sum[8][2] ,
         \ADDER_IN_from_sum[8][1] , \ADDER_IN_from_sum[8][0] ,
         \ADDER_IN_from_sum[7][63] , \ADDER_IN_from_sum[7][62] ,
         \ADDER_IN_from_sum[7][61] , \ADDER_IN_from_sum[7][60] ,
         \ADDER_IN_from_sum[7][59] , \ADDER_IN_from_sum[7][58] ,
         \ADDER_IN_from_sum[7][57] , \ADDER_IN_from_sum[7][56] ,
         \ADDER_IN_from_sum[7][55] , \ADDER_IN_from_sum[7][54] ,
         \ADDER_IN_from_sum[7][53] , \ADDER_IN_from_sum[7][52] ,
         \ADDER_IN_from_sum[7][51] , \ADDER_IN_from_sum[7][50] ,
         \ADDER_IN_from_sum[7][49] , \ADDER_IN_from_sum[7][48] ,
         \ADDER_IN_from_sum[7][47] , \ADDER_IN_from_sum[7][46] ,
         \ADDER_IN_from_sum[7][45] , \ADDER_IN_from_sum[7][44] ,
         \ADDER_IN_from_sum[7][43] , \ADDER_IN_from_sum[7][42] ,
         \ADDER_IN_from_sum[7][41] , \ADDER_IN_from_sum[7][40] ,
         \ADDER_IN_from_sum[7][39] , \ADDER_IN_from_sum[7][38] ,
         \ADDER_IN_from_sum[7][37] , \ADDER_IN_from_sum[7][36] ,
         \ADDER_IN_from_sum[7][35] , \ADDER_IN_from_sum[7][34] ,
         \ADDER_IN_from_sum[7][33] , \ADDER_IN_from_sum[7][32] ,
         \ADDER_IN_from_sum[7][31] , \ADDER_IN_from_sum[7][30] ,
         \ADDER_IN_from_sum[7][29] , \ADDER_IN_from_sum[7][28] ,
         \ADDER_IN_from_sum[7][27] , \ADDER_IN_from_sum[7][26] ,
         \ADDER_IN_from_sum[7][25] , \ADDER_IN_from_sum[7][24] ,
         \ADDER_IN_from_sum[7][23] , \ADDER_IN_from_sum[7][22] ,
         \ADDER_IN_from_sum[7][21] , \ADDER_IN_from_sum[7][20] ,
         \ADDER_IN_from_sum[7][19] , \ADDER_IN_from_sum[7][18] ,
         \ADDER_IN_from_sum[7][17] , \ADDER_IN_from_sum[7][16] ,
         \ADDER_IN_from_sum[7][15] , \ADDER_IN_from_sum[7][14] ,
         \ADDER_IN_from_sum[7][13] , \ADDER_IN_from_sum[7][12] ,
         \ADDER_IN_from_sum[7][11] , \ADDER_IN_from_sum[7][10] ,
         \ADDER_IN_from_sum[7][9] , \ADDER_IN_from_sum[7][8] ,
         \ADDER_IN_from_sum[7][7] , \ADDER_IN_from_sum[7][6] ,
         \ADDER_IN_from_sum[7][5] , \ADDER_IN_from_sum[7][4] ,
         \ADDER_IN_from_sum[7][3] , \ADDER_IN_from_sum[7][2] ,
         \ADDER_IN_from_sum[7][1] , \ADDER_IN_from_sum[7][0] ,
         \ADDER_IN_from_sum[6][63] , \ADDER_IN_from_sum[6][62] ,
         \ADDER_IN_from_sum[6][61] , \ADDER_IN_from_sum[6][60] ,
         \ADDER_IN_from_sum[6][59] , \ADDER_IN_from_sum[6][58] ,
         \ADDER_IN_from_sum[6][57] , \ADDER_IN_from_sum[6][56] ,
         \ADDER_IN_from_sum[6][55] , \ADDER_IN_from_sum[6][54] ,
         \ADDER_IN_from_sum[6][53] , \ADDER_IN_from_sum[6][52] ,
         \ADDER_IN_from_sum[6][51] , \ADDER_IN_from_sum[6][50] ,
         \ADDER_IN_from_sum[6][49] , \ADDER_IN_from_sum[6][48] ,
         \ADDER_IN_from_sum[6][47] , \ADDER_IN_from_sum[6][46] ,
         \ADDER_IN_from_sum[6][45] , \ADDER_IN_from_sum[6][44] ,
         \ADDER_IN_from_sum[6][43] , \ADDER_IN_from_sum[6][42] ,
         \ADDER_IN_from_sum[6][41] , \ADDER_IN_from_sum[6][40] ,
         \ADDER_IN_from_sum[6][39] , \ADDER_IN_from_sum[6][38] ,
         \ADDER_IN_from_sum[6][37] , \ADDER_IN_from_sum[6][36] ,
         \ADDER_IN_from_sum[6][35] , \ADDER_IN_from_sum[6][34] ,
         \ADDER_IN_from_sum[6][33] , \ADDER_IN_from_sum[6][32] ,
         \ADDER_IN_from_sum[6][31] , \ADDER_IN_from_sum[6][30] ,
         \ADDER_IN_from_sum[6][29] , \ADDER_IN_from_sum[6][28] ,
         \ADDER_IN_from_sum[6][27] , \ADDER_IN_from_sum[6][26] ,
         \ADDER_IN_from_sum[6][25] , \ADDER_IN_from_sum[6][24] ,
         \ADDER_IN_from_sum[6][23] , \ADDER_IN_from_sum[6][22] ,
         \ADDER_IN_from_sum[6][21] , \ADDER_IN_from_sum[6][20] ,
         \ADDER_IN_from_sum[6][19] , \ADDER_IN_from_sum[6][18] ,
         \ADDER_IN_from_sum[6][17] , \ADDER_IN_from_sum[6][16] ,
         \ADDER_IN_from_sum[6][15] , \ADDER_IN_from_sum[6][14] ,
         \ADDER_IN_from_sum[6][13] , \ADDER_IN_from_sum[6][12] ,
         \ADDER_IN_from_sum[6][11] , \ADDER_IN_from_sum[6][10] ,
         \ADDER_IN_from_sum[6][9] , \ADDER_IN_from_sum[6][8] ,
         \ADDER_IN_from_sum[6][7] , \ADDER_IN_from_sum[6][6] ,
         \ADDER_IN_from_sum[6][5] , \ADDER_IN_from_sum[6][4] ,
         \ADDER_IN_from_sum[6][3] , \ADDER_IN_from_sum[6][2] ,
         \ADDER_IN_from_sum[6][1] , \ADDER_IN_from_sum[6][0] ,
         \ADDER_IN_from_sum[5][63] , \ADDER_IN_from_sum[5][62] ,
         \ADDER_IN_from_sum[5][61] , \ADDER_IN_from_sum[5][60] ,
         \ADDER_IN_from_sum[5][59] , \ADDER_IN_from_sum[5][58] ,
         \ADDER_IN_from_sum[5][57] , \ADDER_IN_from_sum[5][56] ,
         \ADDER_IN_from_sum[5][55] , \ADDER_IN_from_sum[5][54] ,
         \ADDER_IN_from_sum[5][53] , \ADDER_IN_from_sum[5][52] ,
         \ADDER_IN_from_sum[5][51] , \ADDER_IN_from_sum[5][50] ,
         \ADDER_IN_from_sum[5][49] , \ADDER_IN_from_sum[5][48] ,
         \ADDER_IN_from_sum[5][47] , \ADDER_IN_from_sum[5][46] ,
         \ADDER_IN_from_sum[5][45] , \ADDER_IN_from_sum[5][44] ,
         \ADDER_IN_from_sum[5][43] , \ADDER_IN_from_sum[5][42] ,
         \ADDER_IN_from_sum[5][41] , \ADDER_IN_from_sum[5][40] ,
         \ADDER_IN_from_sum[5][39] , \ADDER_IN_from_sum[5][38] ,
         \ADDER_IN_from_sum[5][37] , \ADDER_IN_from_sum[5][36] ,
         \ADDER_IN_from_sum[5][35] , \ADDER_IN_from_sum[5][34] ,
         \ADDER_IN_from_sum[5][33] , \ADDER_IN_from_sum[5][32] ,
         \ADDER_IN_from_sum[5][31] , \ADDER_IN_from_sum[5][30] ,
         \ADDER_IN_from_sum[5][29] , \ADDER_IN_from_sum[5][28] ,
         \ADDER_IN_from_sum[5][27] , \ADDER_IN_from_sum[5][26] ,
         \ADDER_IN_from_sum[5][25] , \ADDER_IN_from_sum[5][24] ,
         \ADDER_IN_from_sum[5][23] , \ADDER_IN_from_sum[5][22] ,
         \ADDER_IN_from_sum[5][21] , \ADDER_IN_from_sum[5][20] ,
         \ADDER_IN_from_sum[5][19] , \ADDER_IN_from_sum[5][18] ,
         \ADDER_IN_from_sum[5][17] , \ADDER_IN_from_sum[5][16] ,
         \ADDER_IN_from_sum[5][15] , \ADDER_IN_from_sum[5][14] ,
         \ADDER_IN_from_sum[5][13] , \ADDER_IN_from_sum[5][12] ,
         \ADDER_IN_from_sum[5][11] , \ADDER_IN_from_sum[5][10] ,
         \ADDER_IN_from_sum[5][9] , \ADDER_IN_from_sum[5][8] ,
         \ADDER_IN_from_sum[5][7] , \ADDER_IN_from_sum[5][6] ,
         \ADDER_IN_from_sum[5][5] , \ADDER_IN_from_sum[5][4] ,
         \ADDER_IN_from_sum[5][3] , \ADDER_IN_from_sum[5][2] ,
         \ADDER_IN_from_sum[5][1] , \ADDER_IN_from_sum[5][0] ,
         \ADDER_IN_from_sum[4][63] , \ADDER_IN_from_sum[4][62] ,
         \ADDER_IN_from_sum[4][61] , \ADDER_IN_from_sum[4][60] ,
         \ADDER_IN_from_sum[4][59] , \ADDER_IN_from_sum[4][58] ,
         \ADDER_IN_from_sum[4][57] , \ADDER_IN_from_sum[4][56] ,
         \ADDER_IN_from_sum[4][55] , \ADDER_IN_from_sum[4][54] ,
         \ADDER_IN_from_sum[4][53] , \ADDER_IN_from_sum[4][52] ,
         \ADDER_IN_from_sum[4][51] , \ADDER_IN_from_sum[4][50] ,
         \ADDER_IN_from_sum[4][49] , \ADDER_IN_from_sum[4][48] ,
         \ADDER_IN_from_sum[4][47] , \ADDER_IN_from_sum[4][46] ,
         \ADDER_IN_from_sum[4][45] , \ADDER_IN_from_sum[4][44] ,
         \ADDER_IN_from_sum[4][43] , \ADDER_IN_from_sum[4][42] ,
         \ADDER_IN_from_sum[4][41] , \ADDER_IN_from_sum[4][40] ,
         \ADDER_IN_from_sum[4][39] , \ADDER_IN_from_sum[4][38] ,
         \ADDER_IN_from_sum[4][37] , \ADDER_IN_from_sum[4][36] ,
         \ADDER_IN_from_sum[4][35] , \ADDER_IN_from_sum[4][34] ,
         \ADDER_IN_from_sum[4][33] , \ADDER_IN_from_sum[4][32] ,
         \ADDER_IN_from_sum[4][31] , \ADDER_IN_from_sum[4][30] ,
         \ADDER_IN_from_sum[4][29] , \ADDER_IN_from_sum[4][28] ,
         \ADDER_IN_from_sum[4][27] , \ADDER_IN_from_sum[4][26] ,
         \ADDER_IN_from_sum[4][25] , \ADDER_IN_from_sum[4][24] ,
         \ADDER_IN_from_sum[4][23] , \ADDER_IN_from_sum[4][22] ,
         \ADDER_IN_from_sum[4][21] , \ADDER_IN_from_sum[4][20] ,
         \ADDER_IN_from_sum[4][19] , \ADDER_IN_from_sum[4][18] ,
         \ADDER_IN_from_sum[4][17] , \ADDER_IN_from_sum[4][16] ,
         \ADDER_IN_from_sum[4][15] , \ADDER_IN_from_sum[4][14] ,
         \ADDER_IN_from_sum[4][13] , \ADDER_IN_from_sum[4][12] ,
         \ADDER_IN_from_sum[4][11] , \ADDER_IN_from_sum[4][10] ,
         \ADDER_IN_from_sum[4][9] , \ADDER_IN_from_sum[4][8] ,
         \ADDER_IN_from_sum[4][7] , \ADDER_IN_from_sum[4][6] ,
         \ADDER_IN_from_sum[4][5] , \ADDER_IN_from_sum[4][4] ,
         \ADDER_IN_from_sum[4][3] , \ADDER_IN_from_sum[4][2] ,
         \ADDER_IN_from_sum[4][1] , \ADDER_IN_from_sum[4][0] ,
         \ADDER_IN_from_sum[3][63] , \ADDER_IN_from_sum[3][62] ,
         \ADDER_IN_from_sum[3][61] , \ADDER_IN_from_sum[3][60] ,
         \ADDER_IN_from_sum[3][59] , \ADDER_IN_from_sum[3][58] ,
         \ADDER_IN_from_sum[3][57] , \ADDER_IN_from_sum[3][56] ,
         \ADDER_IN_from_sum[3][55] , \ADDER_IN_from_sum[3][54] ,
         \ADDER_IN_from_sum[3][53] , \ADDER_IN_from_sum[3][52] ,
         \ADDER_IN_from_sum[3][51] , \ADDER_IN_from_sum[3][50] ,
         \ADDER_IN_from_sum[3][49] , \ADDER_IN_from_sum[3][48] ,
         \ADDER_IN_from_sum[3][47] , \ADDER_IN_from_sum[3][46] ,
         \ADDER_IN_from_sum[3][45] , \ADDER_IN_from_sum[3][44] ,
         \ADDER_IN_from_sum[3][43] , \ADDER_IN_from_sum[3][42] ,
         \ADDER_IN_from_sum[3][41] , \ADDER_IN_from_sum[3][40] ,
         \ADDER_IN_from_sum[3][39] , \ADDER_IN_from_sum[3][38] ,
         \ADDER_IN_from_sum[3][37] , \ADDER_IN_from_sum[3][36] ,
         \ADDER_IN_from_sum[3][35] , \ADDER_IN_from_sum[3][34] ,
         \ADDER_IN_from_sum[3][33] , \ADDER_IN_from_sum[3][32] ,
         \ADDER_IN_from_sum[3][31] , \ADDER_IN_from_sum[3][30] ,
         \ADDER_IN_from_sum[3][29] , \ADDER_IN_from_sum[3][28] ,
         \ADDER_IN_from_sum[3][27] , \ADDER_IN_from_sum[3][26] ,
         \ADDER_IN_from_sum[3][25] , \ADDER_IN_from_sum[3][24] ,
         \ADDER_IN_from_sum[3][23] , \ADDER_IN_from_sum[3][22] ,
         \ADDER_IN_from_sum[3][21] , \ADDER_IN_from_sum[3][20] ,
         \ADDER_IN_from_sum[3][19] , \ADDER_IN_from_sum[3][18] ,
         \ADDER_IN_from_sum[3][17] , \ADDER_IN_from_sum[3][16] ,
         \ADDER_IN_from_sum[3][15] , \ADDER_IN_from_sum[3][14] ,
         \ADDER_IN_from_sum[3][13] , \ADDER_IN_from_sum[3][12] ,
         \ADDER_IN_from_sum[3][11] , \ADDER_IN_from_sum[3][10] ,
         \ADDER_IN_from_sum[3][9] , \ADDER_IN_from_sum[3][8] ,
         \ADDER_IN_from_sum[3][7] , \ADDER_IN_from_sum[3][6] ,
         \ADDER_IN_from_sum[3][5] , \ADDER_IN_from_sum[3][4] ,
         \ADDER_IN_from_sum[3][3] , \ADDER_IN_from_sum[3][2] ,
         \ADDER_IN_from_sum[3][1] , \ADDER_IN_from_sum[3][0] ,
         \ADDER_IN_from_sum[2][63] , \ADDER_IN_from_sum[2][62] ,
         \ADDER_IN_from_sum[2][61] , \ADDER_IN_from_sum[2][60] ,
         \ADDER_IN_from_sum[2][59] , \ADDER_IN_from_sum[2][58] ,
         \ADDER_IN_from_sum[2][57] , \ADDER_IN_from_sum[2][56] ,
         \ADDER_IN_from_sum[2][55] , \ADDER_IN_from_sum[2][54] ,
         \ADDER_IN_from_sum[2][53] , \ADDER_IN_from_sum[2][52] ,
         \ADDER_IN_from_sum[2][51] , \ADDER_IN_from_sum[2][50] ,
         \ADDER_IN_from_sum[2][49] , \ADDER_IN_from_sum[2][48] ,
         \ADDER_IN_from_sum[2][47] , \ADDER_IN_from_sum[2][46] ,
         \ADDER_IN_from_sum[2][45] , \ADDER_IN_from_sum[2][44] ,
         \ADDER_IN_from_sum[2][43] , \ADDER_IN_from_sum[2][42] ,
         \ADDER_IN_from_sum[2][41] , \ADDER_IN_from_sum[2][40] ,
         \ADDER_IN_from_sum[2][39] , \ADDER_IN_from_sum[2][38] ,
         \ADDER_IN_from_sum[2][37] , \ADDER_IN_from_sum[2][36] ,
         \ADDER_IN_from_sum[2][35] , \ADDER_IN_from_sum[2][34] ,
         \ADDER_IN_from_sum[2][33] , \ADDER_IN_from_sum[2][32] ,
         \ADDER_IN_from_sum[2][31] , \ADDER_IN_from_sum[2][30] ,
         \ADDER_IN_from_sum[2][29] , \ADDER_IN_from_sum[2][28] ,
         \ADDER_IN_from_sum[2][27] , \ADDER_IN_from_sum[2][26] ,
         \ADDER_IN_from_sum[2][25] , \ADDER_IN_from_sum[2][24] ,
         \ADDER_IN_from_sum[2][23] , \ADDER_IN_from_sum[2][22] ,
         \ADDER_IN_from_sum[2][21] , \ADDER_IN_from_sum[2][20] ,
         \ADDER_IN_from_sum[2][19] , \ADDER_IN_from_sum[2][18] ,
         \ADDER_IN_from_sum[2][17] , \ADDER_IN_from_sum[2][16] ,
         \ADDER_IN_from_sum[2][15] , \ADDER_IN_from_sum[2][14] ,
         \ADDER_IN_from_sum[2][13] , \ADDER_IN_from_sum[2][12] ,
         \ADDER_IN_from_sum[2][11] , \ADDER_IN_from_sum[2][10] ,
         \ADDER_IN_from_sum[2][9] , \ADDER_IN_from_sum[2][8] ,
         \ADDER_IN_from_sum[2][7] , \ADDER_IN_from_sum[2][6] ,
         \ADDER_IN_from_sum[2][5] , \ADDER_IN_from_sum[2][4] ,
         \ADDER_IN_from_sum[2][3] , \ADDER_IN_from_sum[2][2] ,
         \ADDER_IN_from_sum[2][1] , \ADDER_IN_from_sum[2][0] ,
         \ADDER_IN_from_sum[1][63] , \ADDER_IN_from_sum[1][62] ,
         \ADDER_IN_from_sum[1][61] , \ADDER_IN_from_sum[1][60] ,
         \ADDER_IN_from_sum[1][59] , \ADDER_IN_from_sum[1][58] ,
         \ADDER_IN_from_sum[1][57] , \ADDER_IN_from_sum[1][56] ,
         \ADDER_IN_from_sum[1][55] , \ADDER_IN_from_sum[1][54] ,
         \ADDER_IN_from_sum[1][53] , \ADDER_IN_from_sum[1][52] ,
         \ADDER_IN_from_sum[1][51] , \ADDER_IN_from_sum[1][50] ,
         \ADDER_IN_from_sum[1][49] , \ADDER_IN_from_sum[1][48] ,
         \ADDER_IN_from_sum[1][47] , \ADDER_IN_from_sum[1][46] ,
         \ADDER_IN_from_sum[1][45] , \ADDER_IN_from_sum[1][44] ,
         \ADDER_IN_from_sum[1][43] , \ADDER_IN_from_sum[1][42] ,
         \ADDER_IN_from_sum[1][41] , \ADDER_IN_from_sum[1][40] ,
         \ADDER_IN_from_sum[1][39] , \ADDER_IN_from_sum[1][38] ,
         \ADDER_IN_from_sum[1][37] , \ADDER_IN_from_sum[1][36] ,
         \ADDER_IN_from_sum[1][35] , \ADDER_IN_from_sum[1][34] ,
         \ADDER_IN_from_sum[1][33] , \ADDER_IN_from_sum[1][32] ,
         \ADDER_IN_from_sum[1][31] , \ADDER_IN_from_sum[1][30] ,
         \ADDER_IN_from_sum[1][29] , \ADDER_IN_from_sum[1][28] ,
         \ADDER_IN_from_sum[1][27] , \ADDER_IN_from_sum[1][26] ,
         \ADDER_IN_from_sum[1][25] , \ADDER_IN_from_sum[1][24] ,
         \ADDER_IN_from_sum[1][23] , \ADDER_IN_from_sum[1][22] ,
         \ADDER_IN_from_sum[1][21] , \ADDER_IN_from_sum[1][20] ,
         \ADDER_IN_from_sum[1][19] , \ADDER_IN_from_sum[1][18] ,
         \ADDER_IN_from_sum[1][17] , \ADDER_IN_from_sum[1][16] ,
         \ADDER_IN_from_sum[1][15] , \ADDER_IN_from_sum[1][14] ,
         \ADDER_IN_from_sum[1][13] , \ADDER_IN_from_sum[1][12] ,
         \ADDER_IN_from_sum[1][11] , \ADDER_IN_from_sum[1][10] ,
         \ADDER_IN_from_sum[1][9] , \ADDER_IN_from_sum[1][8] ,
         \ADDER_IN_from_sum[1][7] , \ADDER_IN_from_sum[1][6] ,
         \ADDER_IN_from_sum[1][5] , \ADDER_IN_from_sum[1][4] ,
         \ADDER_IN_from_sum[1][3] , \ADDER_IN_from_sum[1][2] ,
         \ADDER_IN_from_sum[1][1] , \ADDER_IN_from_sum[1][0] ,
         \ADDER_IN_from_sum[0][63] , \ADDER_IN_from_sum[0][62] ,
         \ADDER_IN_from_sum[0][61] , \ADDER_IN_from_sum[0][60] ,
         \ADDER_IN_from_sum[0][59] , \ADDER_IN_from_sum[0][58] ,
         \ADDER_IN_from_sum[0][57] , \ADDER_IN_from_sum[0][56] ,
         \ADDER_IN_from_sum[0][55] , \ADDER_IN_from_sum[0][54] ,
         \ADDER_IN_from_sum[0][53] , \ADDER_IN_from_sum[0][52] ,
         \ADDER_IN_from_sum[0][51] , \ADDER_IN_from_sum[0][50] ,
         \ADDER_IN_from_sum[0][49] , \ADDER_IN_from_sum[0][48] ,
         \ADDER_IN_from_sum[0][47] , \ADDER_IN_from_sum[0][46] ,
         \ADDER_IN_from_sum[0][45] , \ADDER_IN_from_sum[0][44] ,
         \ADDER_IN_from_sum[0][43] , \ADDER_IN_from_sum[0][42] ,
         \ADDER_IN_from_sum[0][41] , \ADDER_IN_from_sum[0][40] ,
         \ADDER_IN_from_sum[0][39] , \ADDER_IN_from_sum[0][38] ,
         \ADDER_IN_from_sum[0][37] , \ADDER_IN_from_sum[0][36] ,
         \ADDER_IN_from_sum[0][35] , \ADDER_IN_from_sum[0][34] ,
         \ADDER_IN_from_sum[0][33] , \ADDER_IN_from_sum[0][32] ,
         \ADDER_IN_from_sum[0][31] , \ADDER_IN_from_sum[0][30] ,
         \ADDER_IN_from_sum[0][29] , \ADDER_IN_from_sum[0][28] ,
         \ADDER_IN_from_sum[0][27] , \ADDER_IN_from_sum[0][26] ,
         \ADDER_IN_from_sum[0][25] , \ADDER_IN_from_sum[0][24] ,
         \ADDER_IN_from_sum[0][23] , \ADDER_IN_from_sum[0][22] ,
         \ADDER_IN_from_sum[0][21] , \ADDER_IN_from_sum[0][20] ,
         \ADDER_IN_from_sum[0][19] , \ADDER_IN_from_sum[0][18] ,
         \ADDER_IN_from_sum[0][17] , \ADDER_IN_from_sum[0][16] ,
         \ADDER_IN_from_sum[0][15] , \ADDER_IN_from_sum[0][14] ,
         \ADDER_IN_from_sum[0][13] , \ADDER_IN_from_sum[0][12] ,
         \ADDER_IN_from_sum[0][11] , \ADDER_IN_from_sum[0][10] ,
         \ADDER_IN_from_sum[0][9] , \ADDER_IN_from_sum[0][8] ,
         \ADDER_IN_from_sum[0][7] , \ADDER_IN_from_sum[0][6] ,
         \ADDER_IN_from_sum[0][5] , \ADDER_IN_from_sum[0][4] ,
         \ADDER_IN_from_sum[0][3] , \ADDER_IN_from_sum[0][2] ,
         \ADDER_IN_from_sum[0][1] , \ADDER_IN_from_sum[0][0] , n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691;
  wire   [31:0] in_1;
  wire   [31:0] in_2;
  wire   [47:0] Encoder_out;

  FD_GENERIC_NBIT32_0 reg_1 ( .D(INPUT_1), .CLK(Clk), .RESET(reset), .Q(in_1)
         );
  FD_GENERIC_NBIT32_1 reg_2 ( .D(INPUT_2), .CLK(Clk), .RESET(reset), .Q(in_2)
         );
  complement_NBIT64_0 complement_A_signal_0 ( .A({n673, n674, n648, n641, n674, 
        n655, n649, n643, n674, n655, n649, n644, n674, n655, n649, n643, n674, 
        n655, n649, n644, n674, n655, n648, n644, n674, n653, n674, n655, n653, 
        n674, n648, n644, n674, n627, n623, n617, n616, n612, n609, n604, n601, 
        n597, n593, n586, n583, n575, n572, n566, n562, n555, n554, n550, n546, 
        n540, n539, n536, n533, in_1[6], n525, n496, n494, n516, in_1[1], n497}), .Y({\negative_inputs[0][63] , \negative_inputs[0][62] , 
        \negative_inputs[0][61] , \negative_inputs[0][60] , 
        \negative_inputs[0][59] , \negative_inputs[0][58] , 
        \negative_inputs[0][57] , \negative_inputs[0][56] , 
        \negative_inputs[0][55] , \negative_inputs[0][54] , 
        \negative_inputs[0][53] , \negative_inputs[0][52] , 
        \negative_inputs[0][51] , \negative_inputs[0][50] , 
        \negative_inputs[0][49] , \negative_inputs[0][48] , 
        \negative_inputs[0][47] , \negative_inputs[0][46] , 
        \negative_inputs[0][45] , \negative_inputs[0][44] , 
        \negative_inputs[0][43] , \negative_inputs[0][42] , 
        \negative_inputs[0][41] , \negative_inputs[0][40] , 
        \negative_inputs[0][39] , \negative_inputs[0][38] , 
        \negative_inputs[0][37] , \negative_inputs[0][36] , 
        \negative_inputs[0][35] , \negative_inputs[0][34] , 
        \negative_inputs[0][33] , \negative_inputs[0][32] , 
        \negative_inputs[0][31] , \negative_inputs[0][30] , 
        \negative_inputs[0][29] , \negative_inputs[0][28] , 
        \negative_inputs[0][27] , \negative_inputs[0][26] , 
        \negative_inputs[0][25] , \negative_inputs[0][24] , 
        \negative_inputs[0][23] , \negative_inputs[0][22] , 
        \negative_inputs[0][21] , \negative_inputs[0][20] , 
        \negative_inputs[0][19] , \negative_inputs[0][18] , 
        \negative_inputs[0][17] , \negative_inputs[0][16] , 
        \negative_inputs[0][15] , \negative_inputs[0][14] , 
        \negative_inputs[0][13] , \negative_inputs[0][12] , 
        \negative_inputs[0][11] , \negative_inputs[0][10] , 
        \negative_inputs[0][9] , \negative_inputs[0][8] , 
        \negative_inputs[0][7] , \negative_inputs[0][6] , 
        \negative_inputs[0][5] , \negative_inputs[0][4] , 
        \negative_inputs[0][3] , \negative_inputs[0][2] , 
        \negative_inputs[0][1] , \negative_inputs[0][0] }) );
  complement_NBIT64_31 complement_A_signal_1 ( .A({n656, n673, n654, n674, 
        n673, n673, n673, n673, n673, n673, n673, n673, n673, n673, n674, n674, 
        n674, n674, n674, n674, n674, n674, n674, n673, n657, n652, n673, n673, 
        n657, n674, n674, n674, n628, n625, n619, n616, n613, n610, n607, n601, 
        n598, n595, n589, n583, n576, n573, n567, n564, n557, n553, n551, n545, 
        n542, n539, n536, n533, n529, n528, n506, n520, n516, n512, n509, 1'b0}), .Y({\negative_inputs[1][63] , \negative_inputs[1][62] , 
        \negative_inputs[1][61] , \negative_inputs[1][60] , 
        \negative_inputs[1][59] , \negative_inputs[1][58] , 
        \negative_inputs[1][57] , \negative_inputs[1][56] , 
        \negative_inputs[1][55] , \negative_inputs[1][54] , 
        \negative_inputs[1][53] , \negative_inputs[1][52] , 
        \negative_inputs[1][51] , \negative_inputs[1][50] , 
        \negative_inputs[1][49] , \negative_inputs[1][48] , 
        \negative_inputs[1][47] , \negative_inputs[1][46] , 
        \negative_inputs[1][45] , \negative_inputs[1][44] , 
        \negative_inputs[1][43] , \negative_inputs[1][42] , 
        \negative_inputs[1][41] , \negative_inputs[1][40] , 
        \negative_inputs[1][39] , \negative_inputs[1][38] , 
        \negative_inputs[1][37] , \negative_inputs[1][36] , 
        \negative_inputs[1][35] , \negative_inputs[1][34] , 
        \negative_inputs[1][33] , \negative_inputs[1][32] , 
        \negative_inputs[1][31] , \negative_inputs[1][30] , 
        \negative_inputs[1][29] , \negative_inputs[1][28] , 
        \negative_inputs[1][27] , \negative_inputs[1][26] , 
        \negative_inputs[1][25] , \negative_inputs[1][24] , 
        \negative_inputs[1][23] , \negative_inputs[1][22] , 
        \negative_inputs[1][21] , \negative_inputs[1][20] , 
        \negative_inputs[1][19] , \negative_inputs[1][18] , 
        \negative_inputs[1][17] , \negative_inputs[1][16] , 
        \negative_inputs[1][15] , \negative_inputs[1][14] , 
        \negative_inputs[1][13] , \negative_inputs[1][12] , 
        \negative_inputs[1][11] , \negative_inputs[1][10] , 
        \negative_inputs[1][9] , \negative_inputs[1][8] , 
        \negative_inputs[1][7] , \negative_inputs[1][6] , 
        \negative_inputs[1][5] , \negative_inputs[1][4] , 
        \negative_inputs[1][3] , \negative_inputs[1][2] , 
        \negative_inputs[1][1] , \negative_inputs[1][0] }) );
  complement_NBIT64_30 complement_A_signal_2 ( .A({n673, n674, n648, n643, 
        n674, n655, n648, n643, n674, n656, n648, n643, n674, n656, n648, n643, 
        n674, n655, n648, n642, n674, n653, n674, n654, n653, n674, n648, n642, 
        n674, n653, n674, n627, n623, n617, n616, n612, n609, n604, n601, n597, 
        n593, n586, n583, n575, n571, n567, n562, n555, n554, n550, n546, n540, 
        n537, n535, n531, n529, n526, n505, n519, n502, n512, n508, 1'b0, 1'b0}), .Y({\negative_inputs[2][63] , \negative_inputs[2][62] , 
        \negative_inputs[2][61] , \negative_inputs[2][60] , 
        \negative_inputs[2][59] , \negative_inputs[2][58] , 
        \negative_inputs[2][57] , \negative_inputs[2][56] , 
        \negative_inputs[2][55] , \negative_inputs[2][54] , 
        \negative_inputs[2][53] , \negative_inputs[2][52] , 
        \negative_inputs[2][51] , \negative_inputs[2][50] , 
        \negative_inputs[2][49] , \negative_inputs[2][48] , 
        \negative_inputs[2][47] , \negative_inputs[2][46] , 
        \negative_inputs[2][45] , \negative_inputs[2][44] , 
        \negative_inputs[2][43] , \negative_inputs[2][42] , 
        \negative_inputs[2][41] , \negative_inputs[2][40] , 
        \negative_inputs[2][39] , \negative_inputs[2][38] , 
        \negative_inputs[2][37] , \negative_inputs[2][36] , 
        \negative_inputs[2][35] , \negative_inputs[2][34] , 
        \negative_inputs[2][33] , \negative_inputs[2][32] , 
        \negative_inputs[2][31] , \negative_inputs[2][30] , 
        \negative_inputs[2][29] , \negative_inputs[2][28] , 
        \negative_inputs[2][27] , \negative_inputs[2][26] , 
        \negative_inputs[2][25] , \negative_inputs[2][24] , 
        \negative_inputs[2][23] , \negative_inputs[2][22] , 
        \negative_inputs[2][21] , \negative_inputs[2][20] , 
        \negative_inputs[2][19] , \negative_inputs[2][18] , 
        \negative_inputs[2][17] , \negative_inputs[2][16] , 
        \negative_inputs[2][15] , \negative_inputs[2][14] , 
        \negative_inputs[2][13] , \negative_inputs[2][12] , 
        \negative_inputs[2][11] , \negative_inputs[2][10] , 
        \negative_inputs[2][9] , \negative_inputs[2][8] , 
        \negative_inputs[2][7] , \negative_inputs[2][6] , 
        \negative_inputs[2][5] , \negative_inputs[2][4] , 
        \negative_inputs[2][3] , \negative_inputs[2][2] , 
        \negative_inputs[2][1] , \negative_inputs[2][0] }) );
  complement_NBIT64_29 complement_A_signal_3 ( .A({n673, n674, n649, n642, 
        n674, n655, n649, n642, n673, n654, n649, n642, n674, n654, n649, n642, 
        n673, n655, n649, n641, n673, n655, n649, n641, n673, n653, n674, n655, 
        n654, n674, n626, n622, n619, n615, n612, n608, n607, n600, n597, n592, 
        n589, n581, n575, n570, n567, n562, n557, n553, n550, n545, n542, n539, 
        n536, n532, n529, n528, n505, in_1[3], n502, n512, n510, 1'b0, 1'b0, 
        1'b0}), .Y({\negative_inputs[3][63] , \negative_inputs[3][62] , 
        \negative_inputs[3][61] , \negative_inputs[3][60] , 
        \negative_inputs[3][59] , \negative_inputs[3][58] , 
        \negative_inputs[3][57] , \negative_inputs[3][56] , 
        \negative_inputs[3][55] , \negative_inputs[3][54] , 
        \negative_inputs[3][53] , \negative_inputs[3][52] , 
        \negative_inputs[3][51] , \negative_inputs[3][50] , 
        \negative_inputs[3][49] , \negative_inputs[3][48] , 
        \negative_inputs[3][47] , \negative_inputs[3][46] , 
        \negative_inputs[3][45] , \negative_inputs[3][44] , 
        \negative_inputs[3][43] , \negative_inputs[3][42] , 
        \negative_inputs[3][41] , \negative_inputs[3][40] , 
        \negative_inputs[3][39] , \negative_inputs[3][38] , 
        \negative_inputs[3][37] , \negative_inputs[3][36] , 
        \negative_inputs[3][35] , \negative_inputs[3][34] , 
        \negative_inputs[3][33] , \negative_inputs[3][32] , 
        \negative_inputs[3][31] , \negative_inputs[3][30] , 
        \negative_inputs[3][29] , \negative_inputs[3][28] , 
        \negative_inputs[3][27] , \negative_inputs[3][26] , 
        \negative_inputs[3][25] , \negative_inputs[3][24] , 
        \negative_inputs[3][23] , \negative_inputs[3][22] , 
        \negative_inputs[3][21] , \negative_inputs[3][20] , 
        \negative_inputs[3][19] , \negative_inputs[3][18] , 
        \negative_inputs[3][17] , \negative_inputs[3][16] , 
        \negative_inputs[3][15] , \negative_inputs[3][14] , 
        \negative_inputs[3][13] , \negative_inputs[3][12] , 
        \negative_inputs[3][11] , \negative_inputs[3][10] , 
        \negative_inputs[3][9] , \negative_inputs[3][8] , 
        \negative_inputs[3][7] , \negative_inputs[3][6] , 
        \negative_inputs[3][5] , \negative_inputs[3][4] , 
        \negative_inputs[3][3] , \negative_inputs[3][2] , 
        \negative_inputs[3][1] , \negative_inputs[3][0] }) );
  complement_NBIT64_28 complement_A_signal_4 ( .A({n673, n677, n649, n642, 
        n652, n646, n651, n638, n652, n646, n651, n639, n652, n646, n651, n638, 
        n652, n647, n651, n639, n652, n647, n651, n638, n677, n653, n652, n647, 
        n657, n628, n623, n617, n615, n611, n609, n604, n600, n597, n593, n586, 
        n581, n575, n573, n566, n562, n557, n552, n551, n545, n541, n538, n534, 
        n531, n529, n528, n506, n495, n517, n514, n509, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[4][63] , \negative_inputs[4][62] , 
        \negative_inputs[4][61] , \negative_inputs[4][60] , 
        \negative_inputs[4][59] , \negative_inputs[4][58] , 
        \negative_inputs[4][57] , \negative_inputs[4][56] , 
        \negative_inputs[4][55] , \negative_inputs[4][54] , 
        \negative_inputs[4][53] , \negative_inputs[4][52] , 
        \negative_inputs[4][51] , \negative_inputs[4][50] , 
        \negative_inputs[4][49] , \negative_inputs[4][48] , 
        \negative_inputs[4][47] , \negative_inputs[4][46] , 
        \negative_inputs[4][45] , \negative_inputs[4][44] , 
        \negative_inputs[4][43] , \negative_inputs[4][42] , 
        \negative_inputs[4][41] , \negative_inputs[4][40] , 
        \negative_inputs[4][39] , \negative_inputs[4][38] , 
        \negative_inputs[4][37] , \negative_inputs[4][36] , 
        \negative_inputs[4][35] , \negative_inputs[4][34] , 
        \negative_inputs[4][33] , \negative_inputs[4][32] , 
        \negative_inputs[4][31] , \negative_inputs[4][30] , 
        \negative_inputs[4][29] , \negative_inputs[4][28] , 
        \negative_inputs[4][27] , \negative_inputs[4][26] , 
        \negative_inputs[4][25] , \negative_inputs[4][24] , 
        \negative_inputs[4][23] , \negative_inputs[4][22] , 
        \negative_inputs[4][21] , \negative_inputs[4][20] , 
        \negative_inputs[4][19] , \negative_inputs[4][18] , 
        \negative_inputs[4][17] , \negative_inputs[4][16] , 
        \negative_inputs[4][15] , \negative_inputs[4][14] , 
        \negative_inputs[4][13] , \negative_inputs[4][12] , 
        \negative_inputs[4][11] , \negative_inputs[4][10] , 
        \negative_inputs[4][9] , \negative_inputs[4][8] , 
        \negative_inputs[4][7] , \negative_inputs[4][6] , 
        \negative_inputs[4][5] , \negative_inputs[4][4] , 
        \negative_inputs[4][3] , \negative_inputs[4][2] , 
        \negative_inputs[4][1] , \negative_inputs[4][0] }) );
  complement_NBIT64_27 complement_A_signal_5 ( .A({n673, n677, n647, n641, 
        n677, n655, n647, n642, n677, n654, n648, n641, n677, n654, n648, n641, 
        n677, n654, n647, n641, n677, n654, n647, n642, n677, n654, n677, n655, 
        n627, n625, n618, n614, n613, n609, n605, n599, n598, n593, n587, n580, 
        n576, n571, n566, n564, n556, n554, n549, n545, n541, n538, n534, n531, 
        n529, n528, n506, n499, n518, n513, n509, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[5][63] , \negative_inputs[5][62] , 
        \negative_inputs[5][61] , \negative_inputs[5][60] , 
        \negative_inputs[5][59] , \negative_inputs[5][58] , 
        \negative_inputs[5][57] , \negative_inputs[5][56] , 
        \negative_inputs[5][55] , \negative_inputs[5][54] , 
        \negative_inputs[5][53] , \negative_inputs[5][52] , 
        \negative_inputs[5][51] , \negative_inputs[5][50] , 
        \negative_inputs[5][49] , \negative_inputs[5][48] , 
        \negative_inputs[5][47] , \negative_inputs[5][46] , 
        \negative_inputs[5][45] , \negative_inputs[5][44] , 
        \negative_inputs[5][43] , \negative_inputs[5][42] , 
        \negative_inputs[5][41] , \negative_inputs[5][40] , 
        \negative_inputs[5][39] , \negative_inputs[5][38] , 
        \negative_inputs[5][37] , \negative_inputs[5][36] , 
        \negative_inputs[5][35] , \negative_inputs[5][34] , 
        \negative_inputs[5][33] , \negative_inputs[5][32] , 
        \negative_inputs[5][31] , \negative_inputs[5][30] , 
        \negative_inputs[5][29] , \negative_inputs[5][28] , 
        \negative_inputs[5][27] , \negative_inputs[5][26] , 
        \negative_inputs[5][25] , \negative_inputs[5][24] , 
        \negative_inputs[5][23] , \negative_inputs[5][22] , 
        \negative_inputs[5][21] , \negative_inputs[5][20] , 
        \negative_inputs[5][19] , \negative_inputs[5][18] , 
        \negative_inputs[5][17] , \negative_inputs[5][16] , 
        \negative_inputs[5][15] , \negative_inputs[5][14] , 
        \negative_inputs[5][13] , \negative_inputs[5][12] , 
        \negative_inputs[5][11] , \negative_inputs[5][10] , 
        \negative_inputs[5][9] , \negative_inputs[5][8] , 
        \negative_inputs[5][7] , \negative_inputs[5][6] , 
        \negative_inputs[5][5] , \negative_inputs[5][4] , 
        \negative_inputs[5][3] , \negative_inputs[5][2] , 
        \negative_inputs[5][1] , \negative_inputs[5][0] }) );
  complement_NBIT64_26 complement_A_signal_6 ( .A({n673, n677, n677, n677, 
        n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, 
        n657, n652, n656, n655, n657, n652, n656, n676, n657, n652, n655, n628, 
        n624, n618, n615, n612, n609, n605, n601, n597, n593, n587, n583, n576, 
        n571, n566, n562, n557, n553, n550, n545, n541, n538, n534, n531, n530, 
        n501, n496, n520, n518, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[6][63] , \negative_inputs[6][62] , 
        \negative_inputs[6][61] , \negative_inputs[6][60] , 
        \negative_inputs[6][59] , \negative_inputs[6][58] , 
        \negative_inputs[6][57] , \negative_inputs[6][56] , 
        \negative_inputs[6][55] , \negative_inputs[6][54] , 
        \negative_inputs[6][53] , \negative_inputs[6][52] , 
        \negative_inputs[6][51] , \negative_inputs[6][50] , 
        \negative_inputs[6][49] , \negative_inputs[6][48] , 
        \negative_inputs[6][47] , \negative_inputs[6][46] , 
        \negative_inputs[6][45] , \negative_inputs[6][44] , 
        \negative_inputs[6][43] , \negative_inputs[6][42] , 
        \negative_inputs[6][41] , \negative_inputs[6][40] , 
        \negative_inputs[6][39] , \negative_inputs[6][38] , 
        \negative_inputs[6][37] , \negative_inputs[6][36] , 
        \negative_inputs[6][35] , \negative_inputs[6][34] , 
        \negative_inputs[6][33] , \negative_inputs[6][32] , 
        \negative_inputs[6][31] , \negative_inputs[6][30] , 
        \negative_inputs[6][29] , \negative_inputs[6][28] , 
        \negative_inputs[6][27] , \negative_inputs[6][26] , 
        \negative_inputs[6][25] , \negative_inputs[6][24] , 
        \negative_inputs[6][23] , \negative_inputs[6][22] , 
        \negative_inputs[6][21] , \negative_inputs[6][20] , 
        \negative_inputs[6][19] , \negative_inputs[6][18] , 
        \negative_inputs[6][17] , \negative_inputs[6][16] , 
        \negative_inputs[6][15] , \negative_inputs[6][14] , 
        \negative_inputs[6][13] , \negative_inputs[6][12] , 
        \negative_inputs[6][11] , \negative_inputs[6][10] , 
        \negative_inputs[6][9] , \negative_inputs[6][8] , 
        \negative_inputs[6][7] , \negative_inputs[6][6] , 
        \negative_inputs[6][5] , \negative_inputs[6][4] , 
        \negative_inputs[6][3] , \negative_inputs[6][2] , 
        \negative_inputs[6][1] , \negative_inputs[6][0] }) );
  complement_NBIT64_25 complement_A_signal_7 ( .A({n673, n676, n644, n638, 
        n651, n640, n644, n638, n651, n640, n644, n637, n650, n640, n644, n638, 
        n650, n641, n645, n637, n650, n641, n644, n638, n657, n676, n626, n622, 
        n619, n615, n613, n610, n605, n599, n596, n592, n587, n579, n574, n570, 
        n566, n560, n556, n552, n550, n548, n541, n538, n535, n532, n529, n528, 
        n496, n499, n518, n513, n509, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[7][63] , \negative_inputs[7][62] , 
        \negative_inputs[7][61] , \negative_inputs[7][60] , 
        \negative_inputs[7][59] , \negative_inputs[7][58] , 
        \negative_inputs[7][57] , \negative_inputs[7][56] , 
        \negative_inputs[7][55] , \negative_inputs[7][54] , 
        \negative_inputs[7][53] , \negative_inputs[7][52] , 
        \negative_inputs[7][51] , \negative_inputs[7][50] , 
        \negative_inputs[7][49] , \negative_inputs[7][48] , 
        \negative_inputs[7][47] , \negative_inputs[7][46] , 
        \negative_inputs[7][45] , \negative_inputs[7][44] , 
        \negative_inputs[7][43] , \negative_inputs[7][42] , 
        \negative_inputs[7][41] , \negative_inputs[7][40] , 
        \negative_inputs[7][39] , \negative_inputs[7][38] , 
        \negative_inputs[7][37] , \negative_inputs[7][36] , 
        \negative_inputs[7][35] , \negative_inputs[7][34] , 
        \negative_inputs[7][33] , \negative_inputs[7][32] , 
        \negative_inputs[7][31] , \negative_inputs[7][30] , 
        \negative_inputs[7][29] , \negative_inputs[7][28] , 
        \negative_inputs[7][27] , \negative_inputs[7][26] , 
        \negative_inputs[7][25] , \negative_inputs[7][24] , 
        \negative_inputs[7][23] , \negative_inputs[7][22] , 
        \negative_inputs[7][21] , \negative_inputs[7][20] , 
        \negative_inputs[7][19] , \negative_inputs[7][18] , 
        \negative_inputs[7][17] , \negative_inputs[7][16] , 
        \negative_inputs[7][15] , \negative_inputs[7][14] , 
        \negative_inputs[7][13] , \negative_inputs[7][12] , 
        \negative_inputs[7][11] , \negative_inputs[7][10] , 
        \negative_inputs[7][9] , \negative_inputs[7][8] , 
        \negative_inputs[7][7] , \negative_inputs[7][6] , 
        \negative_inputs[7][5] , \negative_inputs[7][4] , 
        \negative_inputs[7][3] , \negative_inputs[7][2] , 
        \negative_inputs[7][1] , \negative_inputs[7][0] }) );
  complement_NBIT64_24 complement_A_signal_8 ( .A({n673, n676, n647, n643, 
        n645, n637, n650, n639, n645, n637, n650, n640, n644, n638, n649, n640, 
        n644, n638, n649, n640, n644, n636, n650, n640, n676, n627, n623, n617, 
        n615, n613, n609, n604, n600, n597, n593, n586, n581, n575, n571, n565, 
        n561, n555, n553, n549, n548, n541, n538, n535, n532, n529, n528, n496, 
        n494, n503, n515, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[8][63] , \negative_inputs[8][62] , 
        \negative_inputs[8][61] , \negative_inputs[8][60] , 
        \negative_inputs[8][59] , \negative_inputs[8][58] , 
        \negative_inputs[8][57] , \negative_inputs[8][56] , 
        \negative_inputs[8][55] , \negative_inputs[8][54] , 
        \negative_inputs[8][53] , \negative_inputs[8][52] , 
        \negative_inputs[8][51] , \negative_inputs[8][50] , 
        \negative_inputs[8][49] , \negative_inputs[8][48] , 
        \negative_inputs[8][47] , \negative_inputs[8][46] , 
        \negative_inputs[8][45] , \negative_inputs[8][44] , 
        \negative_inputs[8][43] , \negative_inputs[8][42] , 
        \negative_inputs[8][41] , \negative_inputs[8][40] , 
        \negative_inputs[8][39] , \negative_inputs[8][38] , 
        \negative_inputs[8][37] , \negative_inputs[8][36] , 
        \negative_inputs[8][35] , \negative_inputs[8][34] , 
        \negative_inputs[8][33] , \negative_inputs[8][32] , 
        \negative_inputs[8][31] , \negative_inputs[8][30] , 
        \negative_inputs[8][29] , \negative_inputs[8][28] , 
        \negative_inputs[8][27] , \negative_inputs[8][26] , 
        \negative_inputs[8][25] , \negative_inputs[8][24] , 
        \negative_inputs[8][23] , \negative_inputs[8][22] , 
        \negative_inputs[8][21] , \negative_inputs[8][20] , 
        \negative_inputs[8][19] , \negative_inputs[8][18] , 
        \negative_inputs[8][17] , \negative_inputs[8][16] , 
        \negative_inputs[8][15] , \negative_inputs[8][14] , 
        \negative_inputs[8][13] , \negative_inputs[8][12] , 
        \negative_inputs[8][11] , \negative_inputs[8][10] , 
        \negative_inputs[8][9] , \negative_inputs[8][8] , 
        \negative_inputs[8][7] , \negative_inputs[8][6] , 
        \negative_inputs[8][5] , \negative_inputs[8][4] , 
        \negative_inputs[8][3] , \negative_inputs[8][2] , 
        \negative_inputs[8][1] , \negative_inputs[8][0] }) );
  complement_NBIT64_23 complement_A_signal_9 ( .A({n673, n676, n676, n676, 
        n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, 
        n657, n652, n656, n676, n657, n652, n676, n676, n627, n624, n618, n616, 
        n612, n609, n606, n600, n597, n593, n588, n581, n575, n571, n567, n564, 
        n556, n553, n551, n548, n541, n538, n534, n531, n491, n501, n506, n500, 
        n518, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[9][63] , \negative_inputs[9][62] , 
        \negative_inputs[9][61] , \negative_inputs[9][60] , 
        \negative_inputs[9][59] , \negative_inputs[9][58] , 
        \negative_inputs[9][57] , \negative_inputs[9][56] , 
        \negative_inputs[9][55] , \negative_inputs[9][54] , 
        \negative_inputs[9][53] , \negative_inputs[9][52] , 
        \negative_inputs[9][51] , \negative_inputs[9][50] , 
        \negative_inputs[9][49] , \negative_inputs[9][48] , 
        \negative_inputs[9][47] , \negative_inputs[9][46] , 
        \negative_inputs[9][45] , \negative_inputs[9][44] , 
        \negative_inputs[9][43] , \negative_inputs[9][42] , 
        \negative_inputs[9][41] , \negative_inputs[9][40] , 
        \negative_inputs[9][39] , \negative_inputs[9][38] , 
        \negative_inputs[9][37] , \negative_inputs[9][36] , 
        \negative_inputs[9][35] , \negative_inputs[9][34] , 
        \negative_inputs[9][33] , \negative_inputs[9][32] , 
        \negative_inputs[9][31] , \negative_inputs[9][30] , 
        \negative_inputs[9][29] , \negative_inputs[9][28] , 
        \negative_inputs[9][27] , \negative_inputs[9][26] , 
        \negative_inputs[9][25] , \negative_inputs[9][24] , 
        \negative_inputs[9][23] , \negative_inputs[9][22] , 
        \negative_inputs[9][21] , \negative_inputs[9][20] , 
        \negative_inputs[9][19] , \negative_inputs[9][18] , 
        \negative_inputs[9][17] , \negative_inputs[9][16] , 
        \negative_inputs[9][15] , \negative_inputs[9][14] , 
        \negative_inputs[9][13] , \negative_inputs[9][12] , 
        \negative_inputs[9][11] , \negative_inputs[9][10] , 
        \negative_inputs[9][9] , \negative_inputs[9][8] , 
        \negative_inputs[9][7] , \negative_inputs[9][6] , 
        \negative_inputs[9][5] , \negative_inputs[9][4] , 
        \negative_inputs[9][3] , \negative_inputs[9][2] , 
        \negative_inputs[9][1] , \negative_inputs[9][0] }) );
  complement_NBIT64_22 complement_A_signal_10 ( .A({n673, n676, n654, n676, 
        n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, n676, 
        n657, n652, n676, n675, n657, n652, n675, n628, n625, n619, n616, n613, 
        n610, n607, n601, n598, n595, n588, n583, n576, n572, n567, n564, n556, 
        n554, n551, n548, n542, n538, n535, n532, n529, n528, n496, n500, n504, 
        n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[10][63] , \negative_inputs[10][62] , 
        \negative_inputs[10][61] , \negative_inputs[10][60] , 
        \negative_inputs[10][59] , \negative_inputs[10][58] , 
        \negative_inputs[10][57] , \negative_inputs[10][56] , 
        \negative_inputs[10][55] , \negative_inputs[10][54] , 
        \negative_inputs[10][53] , \negative_inputs[10][52] , 
        \negative_inputs[10][51] , \negative_inputs[10][50] , 
        \negative_inputs[10][49] , \negative_inputs[10][48] , 
        \negative_inputs[10][47] , \negative_inputs[10][46] , 
        \negative_inputs[10][45] , \negative_inputs[10][44] , 
        \negative_inputs[10][43] , \negative_inputs[10][42] , 
        \negative_inputs[10][41] , \negative_inputs[10][40] , 
        \negative_inputs[10][39] , \negative_inputs[10][38] , 
        \negative_inputs[10][37] , \negative_inputs[10][36] , 
        \negative_inputs[10][35] , \negative_inputs[10][34] , 
        \negative_inputs[10][33] , \negative_inputs[10][32] , 
        \negative_inputs[10][31] , \negative_inputs[10][30] , 
        \negative_inputs[10][29] , \negative_inputs[10][28] , 
        \negative_inputs[10][27] , \negative_inputs[10][26] , 
        \negative_inputs[10][25] , \negative_inputs[10][24] , 
        \negative_inputs[10][23] , \negative_inputs[10][22] , 
        \negative_inputs[10][21] , \negative_inputs[10][20] , 
        \negative_inputs[10][19] , \negative_inputs[10][18] , 
        \negative_inputs[10][17] , \negative_inputs[10][16] , 
        \negative_inputs[10][15] , \negative_inputs[10][14] , 
        \negative_inputs[10][13] , \negative_inputs[10][12] , 
        \negative_inputs[10][11] , \negative_inputs[10][10] , 
        \negative_inputs[10][9] , \negative_inputs[10][8] , 
        \negative_inputs[10][7] , \negative_inputs[10][6] , 
        \negative_inputs[10][5] , \negative_inputs[10][4] , 
        \negative_inputs[10][3] , \negative_inputs[10][2] , 
        \negative_inputs[10][1] , \negative_inputs[10][0] }) );
  complement_NBIT64_21 complement_A_signal_11 ( .A({n656, n653, n675, n655, 
        n647, n643, n675, n655, n647, n644, n675, n655, n647, n643, n675, n655, 
        n648, n643, n675, n655, n653, n675, n626, n622, n619, n615, n613, n610, 
        n605, n601, n597, n592, n588, n581, n575, n570, n567, n562, n556, n552, 
        n551, n545, n541, n538, n535, n532, n529, n501, n496, n495, n518, n514, 
        n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[11][63] , \negative_inputs[11][62] , 
        \negative_inputs[11][61] , \negative_inputs[11][60] , 
        \negative_inputs[11][59] , \negative_inputs[11][58] , 
        \negative_inputs[11][57] , \negative_inputs[11][56] , 
        \negative_inputs[11][55] , \negative_inputs[11][54] , 
        \negative_inputs[11][53] , \negative_inputs[11][52] , 
        \negative_inputs[11][51] , \negative_inputs[11][50] , 
        \negative_inputs[11][49] , \negative_inputs[11][48] , 
        \negative_inputs[11][47] , \negative_inputs[11][46] , 
        \negative_inputs[11][45] , \negative_inputs[11][44] , 
        \negative_inputs[11][43] , \negative_inputs[11][42] , 
        \negative_inputs[11][41] , \negative_inputs[11][40] , 
        \negative_inputs[11][39] , \negative_inputs[11][38] , 
        \negative_inputs[11][37] , \negative_inputs[11][36] , 
        \negative_inputs[11][35] , \negative_inputs[11][34] , 
        \negative_inputs[11][33] , \negative_inputs[11][32] , 
        \negative_inputs[11][31] , \negative_inputs[11][30] , 
        \negative_inputs[11][29] , \negative_inputs[11][28] , 
        \negative_inputs[11][27] , \negative_inputs[11][26] , 
        \negative_inputs[11][25] , \negative_inputs[11][24] , 
        \negative_inputs[11][23] , \negative_inputs[11][22] , 
        \negative_inputs[11][21] , \negative_inputs[11][20] , 
        \negative_inputs[11][19] , \negative_inputs[11][18] , 
        \negative_inputs[11][17] , \negative_inputs[11][16] , 
        \negative_inputs[11][15] , \negative_inputs[11][14] , 
        \negative_inputs[11][13] , \negative_inputs[11][12] , 
        \negative_inputs[11][11] , \negative_inputs[11][10] , 
        \negative_inputs[11][9] , \negative_inputs[11][8] , 
        \negative_inputs[11][7] , \negative_inputs[11][6] , 
        \negative_inputs[11][5] , \negative_inputs[11][4] , 
        \negative_inputs[11][3] , \negative_inputs[11][2] , 
        \negative_inputs[11][1] , \negative_inputs[11][0] }) );
  complement_NBIT64_20 complement_A_signal_12 ( .A({n657, n652, n675, n653, 
        n656, n675, n654, n657, n675, n636, n654, n675, n675, n636, n654, n675, 
        n675, n636, n654, n675, n675, n626, n625, n617, n616, n611, n610, n604, 
        n601, n596, n595, n588, n583, n574, n571, n567, n564, n555, n554, n549, 
        n548, n540, n538, n535, n532, n530, n528, n506, n500, n504, n515, n507, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[12][63] , \negative_inputs[12][62] , 
        \negative_inputs[12][61] , \negative_inputs[12][60] , 
        \negative_inputs[12][59] , \negative_inputs[12][58] , 
        \negative_inputs[12][57] , \negative_inputs[12][56] , 
        \negative_inputs[12][55] , \negative_inputs[12][54] , 
        \negative_inputs[12][53] , \negative_inputs[12][52] , 
        \negative_inputs[12][51] , \negative_inputs[12][50] , 
        \negative_inputs[12][49] , \negative_inputs[12][48] , 
        \negative_inputs[12][47] , \negative_inputs[12][46] , 
        \negative_inputs[12][45] , \negative_inputs[12][44] , 
        \negative_inputs[12][43] , \negative_inputs[12][42] , 
        \negative_inputs[12][41] , \negative_inputs[12][40] , 
        \negative_inputs[12][39] , \negative_inputs[12][38] , 
        \negative_inputs[12][37] , \negative_inputs[12][36] , 
        \negative_inputs[12][35] , \negative_inputs[12][34] , 
        \negative_inputs[12][33] , \negative_inputs[12][32] , 
        \negative_inputs[12][31] , \negative_inputs[12][30] , 
        \negative_inputs[12][29] , \negative_inputs[12][28] , 
        \negative_inputs[12][27] , \negative_inputs[12][26] , 
        \negative_inputs[12][25] , \negative_inputs[12][24] , 
        \negative_inputs[12][23] , \negative_inputs[12][22] , 
        \negative_inputs[12][21] , \negative_inputs[12][20] , 
        \negative_inputs[12][19] , \negative_inputs[12][18] , 
        \negative_inputs[12][17] , \negative_inputs[12][16] , 
        \negative_inputs[12][15] , \negative_inputs[12][14] , 
        \negative_inputs[12][13] , \negative_inputs[12][12] , 
        \negative_inputs[12][11] , \negative_inputs[12][10] , 
        \negative_inputs[12][9] , \negative_inputs[12][8] , 
        \negative_inputs[12][7] , \negative_inputs[12][6] , 
        \negative_inputs[12][5] , \negative_inputs[12][4] , 
        \negative_inputs[12][3] , \negative_inputs[12][2] , 
        \negative_inputs[12][1] , \negative_inputs[12][0] }) );
  complement_NBIT64_19 complement_A_signal_13 ( .A({n673, n675, n647, n643, 
        n646, n637, n650, n639, n646, n636, n651, n639, n646, n636, n651, n640, 
        n646, n636, n651, n639, n626, n622, n618, n614, n611, n608, n605, n599, 
        n598, n593, n587, n579, n575, n570, n565, n560, n556, n552, n549, n545, 
        n541, n538, n535, n531, n491, n501, n522, n500, n504, n515, n507, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[13][63] , \negative_inputs[13][62] , 
        \negative_inputs[13][61] , \negative_inputs[13][60] , 
        \negative_inputs[13][59] , \negative_inputs[13][58] , 
        \negative_inputs[13][57] , \negative_inputs[13][56] , 
        \negative_inputs[13][55] , \negative_inputs[13][54] , 
        \negative_inputs[13][53] , \negative_inputs[13][52] , 
        \negative_inputs[13][51] , \negative_inputs[13][50] , 
        \negative_inputs[13][49] , \negative_inputs[13][48] , 
        \negative_inputs[13][47] , \negative_inputs[13][46] , 
        \negative_inputs[13][45] , \negative_inputs[13][44] , 
        \negative_inputs[13][43] , \negative_inputs[13][42] , 
        \negative_inputs[13][41] , \negative_inputs[13][40] , 
        \negative_inputs[13][39] , \negative_inputs[13][38] , 
        \negative_inputs[13][37] , \negative_inputs[13][36] , 
        \negative_inputs[13][35] , \negative_inputs[13][34] , 
        \negative_inputs[13][33] , \negative_inputs[13][32] , 
        \negative_inputs[13][31] , \negative_inputs[13][30] , 
        \negative_inputs[13][29] , \negative_inputs[13][28] , 
        \negative_inputs[13][27] , \negative_inputs[13][26] , 
        \negative_inputs[13][25] , \negative_inputs[13][24] , 
        \negative_inputs[13][23] , \negative_inputs[13][22] , 
        \negative_inputs[13][21] , \negative_inputs[13][20] , 
        \negative_inputs[13][19] , \negative_inputs[13][18] , 
        \negative_inputs[13][17] , \negative_inputs[13][16] , 
        \negative_inputs[13][15] , \negative_inputs[13][14] , 
        \negative_inputs[13][13] , \negative_inputs[13][12] , 
        \negative_inputs[13][11] , \negative_inputs[13][10] , 
        \negative_inputs[13][9] , \negative_inputs[13][8] , 
        \negative_inputs[13][7] , \negative_inputs[13][6] , 
        \negative_inputs[13][5] , \negative_inputs[13][4] , 
        \negative_inputs[13][3] , \negative_inputs[13][2] , 
        \negative_inputs[13][1] , \negative_inputs[13][0] }) );
  complement_NBIT64_18 complement_A_signal_14 ( .A({n673, n675, n654, n675, 
        n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, 
        n675, n675, n675, n628, n625, n619, n616, n613, n610, n605, n601, n598, 
        n595, n589, n583, n576, n572, n567, n564, n557, n554, n551, n548, n542, 
        n538, n535, n532, n491, n501, n506, n500, n504, n513, n507, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[14][63] , \negative_inputs[14][62] , 
        \negative_inputs[14][61] , \negative_inputs[14][60] , 
        \negative_inputs[14][59] , \negative_inputs[14][58] , 
        \negative_inputs[14][57] , \negative_inputs[14][56] , 
        \negative_inputs[14][55] , \negative_inputs[14][54] , 
        \negative_inputs[14][53] , \negative_inputs[14][52] , 
        \negative_inputs[14][51] , \negative_inputs[14][50] , 
        \negative_inputs[14][49] , \negative_inputs[14][48] , 
        \negative_inputs[14][47] , \negative_inputs[14][46] , 
        \negative_inputs[14][45] , \negative_inputs[14][44] , 
        \negative_inputs[14][43] , \negative_inputs[14][42] , 
        \negative_inputs[14][41] , \negative_inputs[14][40] , 
        \negative_inputs[14][39] , \negative_inputs[14][38] , 
        \negative_inputs[14][37] , \negative_inputs[14][36] , 
        \negative_inputs[14][35] , \negative_inputs[14][34] , 
        \negative_inputs[14][33] , \negative_inputs[14][32] , 
        \negative_inputs[14][31] , \negative_inputs[14][30] , 
        \negative_inputs[14][29] , \negative_inputs[14][28] , 
        \negative_inputs[14][27] , \negative_inputs[14][26] , 
        \negative_inputs[14][25] , \negative_inputs[14][24] , 
        \negative_inputs[14][23] , \negative_inputs[14][22] , 
        \negative_inputs[14][21] , \negative_inputs[14][20] , 
        \negative_inputs[14][19] , \negative_inputs[14][18] , 
        \negative_inputs[14][17] , \negative_inputs[14][16] , 
        \negative_inputs[14][15] , \negative_inputs[14][14] , 
        \negative_inputs[14][13] , \negative_inputs[14][12] , 
        \negative_inputs[14][11] , \negative_inputs[14][10] , 
        \negative_inputs[14][9] , \negative_inputs[14][8] , 
        \negative_inputs[14][7] , \negative_inputs[14][6] , 
        \negative_inputs[14][5] , \negative_inputs[14][4] , 
        \negative_inputs[14][3] , \negative_inputs[14][2] , 
        \negative_inputs[14][1] , \negative_inputs[14][0] }) );
  complement_NBIT64_17 complement_A_signal_15 ( .A({n673, n675, n675, n675, 
        n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, n675, 
        n657, n652, n628, n624, n618, n615, n613, n610, n607, n600, n598, n595, 
        n587, n581, n575, n573, n567, n564, n557, n554, n550, n548, n542, n538, 
        n534, n532, n491, n528, n496, n500, n504, n514, n507, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[15][63] , \negative_inputs[15][62] , 
        \negative_inputs[15][61] , \negative_inputs[15][60] , 
        \negative_inputs[15][59] , \negative_inputs[15][58] , 
        \negative_inputs[15][57] , \negative_inputs[15][56] , 
        \negative_inputs[15][55] , \negative_inputs[15][54] , 
        \negative_inputs[15][53] , \negative_inputs[15][52] , 
        \negative_inputs[15][51] , \negative_inputs[15][50] , 
        \negative_inputs[15][49] , \negative_inputs[15][48] , 
        \negative_inputs[15][47] , \negative_inputs[15][46] , 
        \negative_inputs[15][45] , \negative_inputs[15][44] , 
        \negative_inputs[15][43] , \negative_inputs[15][42] , 
        \negative_inputs[15][41] , \negative_inputs[15][40] , 
        \negative_inputs[15][39] , \negative_inputs[15][38] , 
        \negative_inputs[15][37] , \negative_inputs[15][36] , 
        \negative_inputs[15][35] , \negative_inputs[15][34] , 
        \negative_inputs[15][33] , \negative_inputs[15][32] , 
        \negative_inputs[15][31] , \negative_inputs[15][30] , 
        \negative_inputs[15][29] , \negative_inputs[15][28] , 
        \negative_inputs[15][27] , \negative_inputs[15][26] , 
        \negative_inputs[15][25] , \negative_inputs[15][24] , 
        \negative_inputs[15][23] , \negative_inputs[15][22] , 
        \negative_inputs[15][21] , \negative_inputs[15][20] , 
        \negative_inputs[15][19] , \negative_inputs[15][18] , 
        \negative_inputs[15][17] , \negative_inputs[15][16] , 
        \negative_inputs[15][15] , \negative_inputs[15][14] , 
        \negative_inputs[15][13] , \negative_inputs[15][12] , 
        \negative_inputs[15][11] , \negative_inputs[15][10] , 
        \negative_inputs[15][9] , \negative_inputs[15][8] , 
        \negative_inputs[15][7] , \negative_inputs[15][6] , 
        \negative_inputs[15][5] , \negative_inputs[15][4] , 
        \negative_inputs[15][3] , \negative_inputs[15][2] , 
        \negative_inputs[15][1] , \negative_inputs[15][0] }) );
  complement_NBIT64_16 complement_A_signal_16 ( .A({n656, n653, n675, n647, 
        n644, n646, n637, n650, n639, n645, n637, n650, n639, n645, n636, n650, 
        n640, n626, n622, n618, n614, n611, n608, n605, n599, n596, n592, n587, 
        n580, n574, n570, n566, n561, n555, n552, n550, n545, n540, n538, n535, 
        n531, n491, n490, n496, n500, n504, n513, n507, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[16][63] , \negative_inputs[16][62] , 
        \negative_inputs[16][61] , \negative_inputs[16][60] , 
        \negative_inputs[16][59] , \negative_inputs[16][58] , 
        \negative_inputs[16][57] , \negative_inputs[16][56] , 
        \negative_inputs[16][55] , \negative_inputs[16][54] , 
        \negative_inputs[16][53] , \negative_inputs[16][52] , 
        \negative_inputs[16][51] , \negative_inputs[16][50] , 
        \negative_inputs[16][49] , \negative_inputs[16][48] , 
        \negative_inputs[16][47] , \negative_inputs[16][46] , 
        \negative_inputs[16][45] , \negative_inputs[16][44] , 
        \negative_inputs[16][43] , \negative_inputs[16][42] , 
        \negative_inputs[16][41] , \negative_inputs[16][40] , 
        \negative_inputs[16][39] , \negative_inputs[16][38] , 
        \negative_inputs[16][37] , \negative_inputs[16][36] , 
        \negative_inputs[16][35] , \negative_inputs[16][34] , 
        \negative_inputs[16][33] , \negative_inputs[16][32] , 
        \negative_inputs[16][31] , \negative_inputs[16][30] , 
        \negative_inputs[16][29] , \negative_inputs[16][28] , 
        \negative_inputs[16][27] , \negative_inputs[16][26] , 
        \negative_inputs[16][25] , \negative_inputs[16][24] , 
        \negative_inputs[16][23] , \negative_inputs[16][22] , 
        \negative_inputs[16][21] , \negative_inputs[16][20] , 
        \negative_inputs[16][19] , \negative_inputs[16][18] , 
        \negative_inputs[16][17] , \negative_inputs[16][16] , 
        \negative_inputs[16][15] , \negative_inputs[16][14] , 
        \negative_inputs[16][13] , \negative_inputs[16][12] , 
        \negative_inputs[16][11] , \negative_inputs[16][10] , 
        \negative_inputs[16][9] , \negative_inputs[16][8] , 
        \negative_inputs[16][7] , \negative_inputs[16][6] , 
        \negative_inputs[16][5] , \negative_inputs[16][4] , 
        \negative_inputs[16][3] , \negative_inputs[16][2] , 
        \negative_inputs[16][1] , \negative_inputs[16][0] }) );
  complement_NBIT64_15 complement_A_signal_17 ( .A({n656, n653, n674, n648, 
        n642, n646, n636, n652, n640, n645, n638, n650, n639, n646, n636, n651, 
        n626, n623, n617, n615, n611, n608, n604, n600, n596, n593, n586, n581, 
        n574, n571, n565, n562, n555, n552, n549, n545, n540, n538, n534, n532, 
        n491, n490, n522, n520, n504, n514, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[17][63] , \negative_inputs[17][62] , 
        \negative_inputs[17][61] , \negative_inputs[17][60] , 
        \negative_inputs[17][59] , \negative_inputs[17][58] , 
        \negative_inputs[17][57] , \negative_inputs[17][56] , 
        \negative_inputs[17][55] , \negative_inputs[17][54] , 
        \negative_inputs[17][53] , \negative_inputs[17][52] , 
        \negative_inputs[17][51] , \negative_inputs[17][50] , 
        \negative_inputs[17][49] , \negative_inputs[17][48] , 
        \negative_inputs[17][47] , \negative_inputs[17][46] , 
        \negative_inputs[17][45] , \negative_inputs[17][44] , 
        \negative_inputs[17][43] , \negative_inputs[17][42] , 
        \negative_inputs[17][41] , \negative_inputs[17][40] , 
        \negative_inputs[17][39] , \negative_inputs[17][38] , 
        \negative_inputs[17][37] , \negative_inputs[17][36] , 
        \negative_inputs[17][35] , \negative_inputs[17][34] , 
        \negative_inputs[17][33] , \negative_inputs[17][32] , 
        \negative_inputs[17][31] , \negative_inputs[17][30] , 
        \negative_inputs[17][29] , \negative_inputs[17][28] , 
        \negative_inputs[17][27] , \negative_inputs[17][26] , 
        \negative_inputs[17][25] , \negative_inputs[17][24] , 
        \negative_inputs[17][23] , \negative_inputs[17][22] , 
        \negative_inputs[17][21] , \negative_inputs[17][20] , 
        \negative_inputs[17][19] , \negative_inputs[17][18] , 
        \negative_inputs[17][17] , \negative_inputs[17][16] , 
        \negative_inputs[17][15] , \negative_inputs[17][14] , 
        \negative_inputs[17][13] , \negative_inputs[17][12] , 
        \negative_inputs[17][11] , \negative_inputs[17][10] , 
        \negative_inputs[17][9] , \negative_inputs[17][8] , 
        \negative_inputs[17][7] , \negative_inputs[17][6] , 
        \negative_inputs[17][5] , \negative_inputs[17][4] , 
        \negative_inputs[17][3] , \negative_inputs[17][2] , 
        \negative_inputs[17][1] , \negative_inputs[17][0] }) );
  complement_NBIT64_14 complement_A_signal_18 ( .A({n656, n654, n674, n649, 
        n643, n646, n636, n650, n639, n646, n637, n650, n639, n652, n646, n627, 
        n622, n618, n614, n612, n608, n605, n599, n597, n592, n587, n579, n575, 
        n570, n565, n560, n556, n552, n549, n545, n541, n538, n535, n532, n491, 
        n490, n522, n499, n504, n513, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[18][63] , \negative_inputs[18][62] , 
        \negative_inputs[18][61] , \negative_inputs[18][60] , 
        \negative_inputs[18][59] , \negative_inputs[18][58] , 
        \negative_inputs[18][57] , \negative_inputs[18][56] , 
        \negative_inputs[18][55] , \negative_inputs[18][54] , 
        \negative_inputs[18][53] , \negative_inputs[18][52] , 
        \negative_inputs[18][51] , \negative_inputs[18][50] , 
        \negative_inputs[18][49] , \negative_inputs[18][48] , 
        \negative_inputs[18][47] , \negative_inputs[18][46] , 
        \negative_inputs[18][45] , \negative_inputs[18][44] , 
        \negative_inputs[18][43] , \negative_inputs[18][42] , 
        \negative_inputs[18][41] , \negative_inputs[18][40] , 
        \negative_inputs[18][39] , \negative_inputs[18][38] , 
        \negative_inputs[18][37] , \negative_inputs[18][36] , 
        \negative_inputs[18][35] , \negative_inputs[18][34] , 
        \negative_inputs[18][33] , \negative_inputs[18][32] , 
        \negative_inputs[18][31] , \negative_inputs[18][30] , 
        \negative_inputs[18][29] , \negative_inputs[18][28] , 
        \negative_inputs[18][27] , \negative_inputs[18][26] , 
        \negative_inputs[18][25] , \negative_inputs[18][24] , 
        \negative_inputs[18][23] , \negative_inputs[18][22] , 
        \negative_inputs[18][21] , \negative_inputs[18][20] , 
        \negative_inputs[18][19] , \negative_inputs[18][18] , 
        \negative_inputs[18][17] , \negative_inputs[18][16] , 
        \negative_inputs[18][15] , \negative_inputs[18][14] , 
        \negative_inputs[18][13] , \negative_inputs[18][12] , 
        \negative_inputs[18][11] , \negative_inputs[18][10] , 
        \negative_inputs[18][9] , \negative_inputs[18][8] , 
        \negative_inputs[18][7] , \negative_inputs[18][6] , 
        \negative_inputs[18][5] , \negative_inputs[18][4] , 
        \negative_inputs[18][3] , \negative_inputs[18][2] , 
        \negative_inputs[18][1] , \negative_inputs[18][0] }) );
  complement_NBIT64_13 complement_A_signal_19 ( .A({n656, n653, n676, n648, 
        n643, n645, n637, n650, n640, n645, n638, n651, n640, n652, n626, n623, 
        n617, n614, n611, n609, n604, n599, n596, n593, n586, n580, n574, n571, 
        n565, n561, n555, n553, n549, n545, n540, n538, n534, n532, n491, n501, 
        n522, n495, n503, n514, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[19][63] , \negative_inputs[19][62] , 
        \negative_inputs[19][61] , \negative_inputs[19][60] , 
        \negative_inputs[19][59] , \negative_inputs[19][58] , 
        \negative_inputs[19][57] , \negative_inputs[19][56] , 
        \negative_inputs[19][55] , \negative_inputs[19][54] , 
        \negative_inputs[19][53] , \negative_inputs[19][52] , 
        \negative_inputs[19][51] , \negative_inputs[19][50] , 
        \negative_inputs[19][49] , \negative_inputs[19][48] , 
        \negative_inputs[19][47] , \negative_inputs[19][46] , 
        \negative_inputs[19][45] , \negative_inputs[19][44] , 
        \negative_inputs[19][43] , \negative_inputs[19][42] , 
        \negative_inputs[19][41] , \negative_inputs[19][40] , 
        \negative_inputs[19][39] , \negative_inputs[19][38] , 
        \negative_inputs[19][37] , \negative_inputs[19][36] , 
        \negative_inputs[19][35] , \negative_inputs[19][34] , 
        \negative_inputs[19][33] , \negative_inputs[19][32] , 
        \negative_inputs[19][31] , \negative_inputs[19][30] , 
        \negative_inputs[19][29] , \negative_inputs[19][28] , 
        \negative_inputs[19][27] , \negative_inputs[19][26] , 
        \negative_inputs[19][25] , \negative_inputs[19][24] , 
        \negative_inputs[19][23] , \negative_inputs[19][22] , 
        \negative_inputs[19][21] , \negative_inputs[19][20] , 
        \negative_inputs[19][19] , \negative_inputs[19][18] , 
        \negative_inputs[19][17] , \negative_inputs[19][16] , 
        \negative_inputs[19][15] , \negative_inputs[19][14] , 
        \negative_inputs[19][13] , \negative_inputs[19][12] , 
        \negative_inputs[19][11] , \negative_inputs[19][10] , 
        \negative_inputs[19][9] , \negative_inputs[19][8] , 
        \negative_inputs[19][7] , \negative_inputs[19][6] , 
        \negative_inputs[19][5] , \negative_inputs[19][4] , 
        \negative_inputs[19][3] , \negative_inputs[19][2] , 
        \negative_inputs[19][1] , \negative_inputs[19][0] }) );
  complement_NBIT64_12 complement_A_signal_20 ( .A({n656, n653, n674, n648, 
        n643, n645, n638, n650, n640, n645, n637, n650, n641, n626, n622, n618, 
        n614, n612, n608, n605, n599, n596, n592, n587, n580, n574, n570, n566, 
        n561, n555, n552, n550, n545, n540, n538, n534, n531, n491, n490, n496, 
        n500, n504, n513, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[20][63] , \negative_inputs[20][62] , 
        \negative_inputs[20][61] , \negative_inputs[20][60] , 
        \negative_inputs[20][59] , \negative_inputs[20][58] , 
        \negative_inputs[20][57] , \negative_inputs[20][56] , 
        \negative_inputs[20][55] , \negative_inputs[20][54] , 
        \negative_inputs[20][53] , \negative_inputs[20][52] , 
        \negative_inputs[20][51] , \negative_inputs[20][50] , 
        \negative_inputs[20][49] , \negative_inputs[20][48] , 
        \negative_inputs[20][47] , \negative_inputs[20][46] , 
        \negative_inputs[20][45] , \negative_inputs[20][44] , 
        \negative_inputs[20][43] , \negative_inputs[20][42] , 
        \negative_inputs[20][41] , \negative_inputs[20][40] , 
        \negative_inputs[20][39] , \negative_inputs[20][38] , 
        \negative_inputs[20][37] , \negative_inputs[20][36] , 
        \negative_inputs[20][35] , \negative_inputs[20][34] , 
        \negative_inputs[20][33] , \negative_inputs[20][32] , 
        \negative_inputs[20][31] , \negative_inputs[20][30] , 
        \negative_inputs[20][29] , \negative_inputs[20][28] , 
        \negative_inputs[20][27] , \negative_inputs[20][26] , 
        \negative_inputs[20][25] , \negative_inputs[20][24] , 
        \negative_inputs[20][23] , \negative_inputs[20][22] , 
        \negative_inputs[20][21] , \negative_inputs[20][20] , 
        \negative_inputs[20][19] , \negative_inputs[20][18] , 
        \negative_inputs[20][17] , \negative_inputs[20][16] , 
        \negative_inputs[20][15] , \negative_inputs[20][14] , 
        \negative_inputs[20][13] , \negative_inputs[20][12] , 
        \negative_inputs[20][11] , \negative_inputs[20][10] , 
        \negative_inputs[20][9] , \negative_inputs[20][8] , 
        \negative_inputs[20][7] , \negative_inputs[20][6] , 
        \negative_inputs[20][5] , \negative_inputs[20][4] , 
        \negative_inputs[20][3] , \negative_inputs[20][2] , 
        \negative_inputs[20][1] , \negative_inputs[20][0] }) );
  complement_NBIT64_11 complement_A_signal_21 ( .A({n656, n653, n674, n649, 
        n642, n644, n637, n651, n640, n645, n638, n650, n626, n623, n617, n615, 
        n611, n609, n605, n600, n596, n592, n586, n581, n574, n571, n565, n562, 
        n555, n552, n549, n545, n540, n538, n535, n532, n491, n490, n522, n520, 
        n504, n514, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[21][63] , \negative_inputs[21][62] , 
        \negative_inputs[21][61] , \negative_inputs[21][60] , 
        \negative_inputs[21][59] , \negative_inputs[21][58] , 
        \negative_inputs[21][57] , \negative_inputs[21][56] , 
        \negative_inputs[21][55] , \negative_inputs[21][54] , 
        \negative_inputs[21][53] , \negative_inputs[21][52] , 
        \negative_inputs[21][51] , \negative_inputs[21][50] , 
        \negative_inputs[21][49] , \negative_inputs[21][48] , 
        \negative_inputs[21][47] , \negative_inputs[21][46] , 
        \negative_inputs[21][45] , \negative_inputs[21][44] , 
        \negative_inputs[21][43] , \negative_inputs[21][42] , 
        \negative_inputs[21][41] , \negative_inputs[21][40] , 
        \negative_inputs[21][39] , \negative_inputs[21][38] , 
        \negative_inputs[21][37] , \negative_inputs[21][36] , 
        \negative_inputs[21][35] , \negative_inputs[21][34] , 
        \negative_inputs[21][33] , \negative_inputs[21][32] , 
        \negative_inputs[21][31] , \negative_inputs[21][30] , 
        \negative_inputs[21][29] , \negative_inputs[21][28] , 
        \negative_inputs[21][27] , \negative_inputs[21][26] , 
        \negative_inputs[21][25] , \negative_inputs[21][24] , 
        \negative_inputs[21][23] , \negative_inputs[21][22] , 
        \negative_inputs[21][21] , \negative_inputs[21][20] , 
        \negative_inputs[21][19] , \negative_inputs[21][18] , 
        \negative_inputs[21][17] , \negative_inputs[21][16] , 
        \negative_inputs[21][15] , \negative_inputs[21][14] , 
        \negative_inputs[21][13] , \negative_inputs[21][12] , 
        \negative_inputs[21][11] , \negative_inputs[21][10] , 
        \negative_inputs[21][9] , \negative_inputs[21][8] , 
        \negative_inputs[21][7] , \negative_inputs[21][6] , 
        \negative_inputs[21][5] , \negative_inputs[21][4] , 
        \negative_inputs[21][3] , \negative_inputs[21][2] , 
        \negative_inputs[21][1] , \negative_inputs[21][0] }) );
  complement_NBIT64_10 complement_A_signal_22 ( .A({n656, n654, n674, n649, 
        n642, n645, n637, n651, n639, n645, n637, n627, n622, n617, n614, n612, 
        n608, n605, n599, n597, n592, n587, n579, n575, n570, n565, n560, n556, 
        n552, n549, n545, n541, n538, n535, n532, n491, n490, n522, n499, n504, 
        n513, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[22][63] , \negative_inputs[22][62] , 
        \negative_inputs[22][61] , \negative_inputs[22][60] , 
        \negative_inputs[22][59] , \negative_inputs[22][58] , 
        \negative_inputs[22][57] , \negative_inputs[22][56] , 
        \negative_inputs[22][55] , \negative_inputs[22][54] , 
        \negative_inputs[22][53] , \negative_inputs[22][52] , 
        \negative_inputs[22][51] , \negative_inputs[22][50] , 
        \negative_inputs[22][49] , \negative_inputs[22][48] , 
        \negative_inputs[22][47] , \negative_inputs[22][46] , 
        \negative_inputs[22][45] , \negative_inputs[22][44] , 
        \negative_inputs[22][43] , \negative_inputs[22][42] , 
        \negative_inputs[22][41] , \negative_inputs[22][40] , 
        \negative_inputs[22][39] , \negative_inputs[22][38] , 
        \negative_inputs[22][37] , \negative_inputs[22][36] , 
        \negative_inputs[22][35] , \negative_inputs[22][34] , 
        \negative_inputs[22][33] , \negative_inputs[22][32] , 
        \negative_inputs[22][31] , \negative_inputs[22][30] , 
        \negative_inputs[22][29] , \negative_inputs[22][28] , 
        \negative_inputs[22][27] , \negative_inputs[22][26] , 
        \negative_inputs[22][25] , \negative_inputs[22][24] , 
        \negative_inputs[22][23] , \negative_inputs[22][22] , 
        \negative_inputs[22][21] , \negative_inputs[22][20] , 
        \negative_inputs[22][19] , \negative_inputs[22][18] , 
        \negative_inputs[22][17] , \negative_inputs[22][16] , 
        \negative_inputs[22][15] , \negative_inputs[22][14] , 
        \negative_inputs[22][13] , \negative_inputs[22][12] , 
        \negative_inputs[22][11] , \negative_inputs[22][10] , 
        \negative_inputs[22][9] , \negative_inputs[22][8] , 
        \negative_inputs[22][7] , \negative_inputs[22][6] , 
        \negative_inputs[22][5] , \negative_inputs[22][4] , 
        \negative_inputs[22][3] , \negative_inputs[22][2] , 
        \negative_inputs[22][1] , \negative_inputs[22][0] }) );
  complement_NBIT64_9 complement_A_signal_23 ( .A({n656, n653, n674, n649, 
        n642, n646, n637, n651, n639, n645, n626, n623, n617, n615, n611, n609, 
        n604, n600, n596, n593, n586, n580, n574, n571, n565, n561, n555, n553, 
        n549, n545, n540, n538, n535, n532, n491, n501, n522, n494, n503, n514, 
        n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[23][63] , \negative_inputs[23][62] , 
        \negative_inputs[23][61] , \negative_inputs[23][60] , 
        \negative_inputs[23][59] , \negative_inputs[23][58] , 
        \negative_inputs[23][57] , \negative_inputs[23][56] , 
        \negative_inputs[23][55] , \negative_inputs[23][54] , 
        \negative_inputs[23][53] , \negative_inputs[23][52] , 
        \negative_inputs[23][51] , \negative_inputs[23][50] , 
        \negative_inputs[23][49] , \negative_inputs[23][48] , 
        \negative_inputs[23][47] , \negative_inputs[23][46] , 
        \negative_inputs[23][45] , \negative_inputs[23][44] , 
        \negative_inputs[23][43] , \negative_inputs[23][42] , 
        \negative_inputs[23][41] , \negative_inputs[23][40] , 
        \negative_inputs[23][39] , \negative_inputs[23][38] , 
        \negative_inputs[23][37] , \negative_inputs[23][36] , 
        \negative_inputs[23][35] , \negative_inputs[23][34] , 
        \negative_inputs[23][33] , \negative_inputs[23][32] , 
        \negative_inputs[23][31] , \negative_inputs[23][30] , 
        \negative_inputs[23][29] , \negative_inputs[23][28] , 
        \negative_inputs[23][27] , \negative_inputs[23][26] , 
        \negative_inputs[23][25] , \negative_inputs[23][24] , 
        \negative_inputs[23][23] , \negative_inputs[23][22] , 
        \negative_inputs[23][21] , \negative_inputs[23][20] , 
        \negative_inputs[23][19] , \negative_inputs[23][18] , 
        \negative_inputs[23][17] , \negative_inputs[23][16] , 
        \negative_inputs[23][15] , \negative_inputs[23][14] , 
        \negative_inputs[23][13] , \negative_inputs[23][12] , 
        \negative_inputs[23][11] , \negative_inputs[23][10] , 
        \negative_inputs[23][9] , \negative_inputs[23][8] , 
        \negative_inputs[23][7] , \negative_inputs[23][6] , 
        \negative_inputs[23][5] , \negative_inputs[23][4] , 
        \negative_inputs[23][3] , \negative_inputs[23][2] , 
        \negative_inputs[23][1] , \negative_inputs[23][0] }) );
  complement_NBIT64_8 complement_A_signal_24 ( .A({n656, n653, n674, n648, 
        n641, n646, n636, n651, n639, n626, n622, n618, n614, n611, n608, n605, 
        n599, n596, n592, n587, n580, n574, n570, n566, n560, n556, n552, n550, 
        n545, n541, n538, n534, n532, n491, n490, n496, n500, n504, n513, n507, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[24][63] , \negative_inputs[24][62] , 
        \negative_inputs[24][61] , \negative_inputs[24][60] , 
        \negative_inputs[24][59] , \negative_inputs[24][58] , 
        \negative_inputs[24][57] , \negative_inputs[24][56] , 
        \negative_inputs[24][55] , \negative_inputs[24][54] , 
        \negative_inputs[24][53] , \negative_inputs[24][52] , 
        \negative_inputs[24][51] , \negative_inputs[24][50] , 
        \negative_inputs[24][49] , \negative_inputs[24][48] , 
        \negative_inputs[24][47] , \negative_inputs[24][46] , 
        \negative_inputs[24][45] , \negative_inputs[24][44] , 
        \negative_inputs[24][43] , \negative_inputs[24][42] , 
        \negative_inputs[24][41] , \negative_inputs[24][40] , 
        \negative_inputs[24][39] , \negative_inputs[24][38] , 
        \negative_inputs[24][37] , \negative_inputs[24][36] , 
        \negative_inputs[24][35] , \negative_inputs[24][34] , 
        \negative_inputs[24][33] , \negative_inputs[24][32] , 
        \negative_inputs[24][31] , \negative_inputs[24][30] , 
        \negative_inputs[24][29] , \negative_inputs[24][28] , 
        \negative_inputs[24][27] , \negative_inputs[24][26] , 
        \negative_inputs[24][25] , \negative_inputs[24][24] , 
        \negative_inputs[24][23] , \negative_inputs[24][22] , 
        \negative_inputs[24][21] , \negative_inputs[24][20] , 
        \negative_inputs[24][19] , \negative_inputs[24][18] , 
        \negative_inputs[24][17] , \negative_inputs[24][16] , 
        \negative_inputs[24][15] , \negative_inputs[24][14] , 
        \negative_inputs[24][13] , \negative_inputs[24][12] , 
        \negative_inputs[24][11] , \negative_inputs[24][10] , 
        \negative_inputs[24][9] , \negative_inputs[24][8] , 
        \negative_inputs[24][7] , \negative_inputs[24][6] , 
        \negative_inputs[24][5] , \negative_inputs[24][4] , 
        \negative_inputs[24][3] , \negative_inputs[24][2] , 
        \negative_inputs[24][1] , \negative_inputs[24][0] }) );
  complement_NBIT64_7 complement_A_signal_25 ( .A({n656, n653, n674, n648, 
        n641, n646, n636, n651, n626, n623, n617, n615, n611, n608, n604, n600, 
        n596, n593, n586, n581, n574, n571, n565, n562, n555, n553, n549, n545, 
        n540, n538, n535, n531, n491, n501, n522, n494, n504, n514, n493, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[25][63] , \negative_inputs[25][62] , 
        \negative_inputs[25][61] , \negative_inputs[25][60] , 
        \negative_inputs[25][59] , \negative_inputs[25][58] , 
        \negative_inputs[25][57] , \negative_inputs[25][56] , 
        \negative_inputs[25][55] , \negative_inputs[25][54] , 
        \negative_inputs[25][53] , \negative_inputs[25][52] , 
        \negative_inputs[25][51] , \negative_inputs[25][50] , 
        \negative_inputs[25][49] , \negative_inputs[25][48] , 
        \negative_inputs[25][47] , \negative_inputs[25][46] , 
        \negative_inputs[25][45] , \negative_inputs[25][44] , 
        \negative_inputs[25][43] , \negative_inputs[25][42] , 
        \negative_inputs[25][41] , \negative_inputs[25][40] , 
        \negative_inputs[25][39] , \negative_inputs[25][38] , 
        \negative_inputs[25][37] , \negative_inputs[25][36] , 
        \negative_inputs[25][35] , \negative_inputs[25][34] , 
        \negative_inputs[25][33] , \negative_inputs[25][32] , 
        \negative_inputs[25][31] , \negative_inputs[25][30] , 
        \negative_inputs[25][29] , \negative_inputs[25][28] , 
        \negative_inputs[25][27] , \negative_inputs[25][26] , 
        \negative_inputs[25][25] , \negative_inputs[25][24] , 
        \negative_inputs[25][23] , \negative_inputs[25][22] , 
        \negative_inputs[25][21] , \negative_inputs[25][20] , 
        \negative_inputs[25][19] , \negative_inputs[25][18] , 
        \negative_inputs[25][17] , \negative_inputs[25][16] , 
        \negative_inputs[25][15] , \negative_inputs[25][14] , 
        \negative_inputs[25][13] , \negative_inputs[25][12] , 
        \negative_inputs[25][11] , \negative_inputs[25][10] , 
        \negative_inputs[25][9] , \negative_inputs[25][8] , 
        \negative_inputs[25][7] , \negative_inputs[25][6] , 
        \negative_inputs[25][5] , \negative_inputs[25][4] , 
        \negative_inputs[25][3] , \negative_inputs[25][2] , 
        \negative_inputs[25][1] , \negative_inputs[25][0] }) );
  complement_NBIT64_6 complement_A_signal_26 ( .A({n656, n653, n674, n647, 
        n642, n645, n638, n627, n622, n618, n614, n612, n608, n605, n599, n597, 
        n592, n587, n579, n575, n570, n566, n560, n556, n552, n550, n545, n541, 
        n538, n534, n532, n530, n490, n522, n499, n504, n513, n507, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[26][63] , \negative_inputs[26][62] , 
        \negative_inputs[26][61] , \negative_inputs[26][60] , 
        \negative_inputs[26][59] , \negative_inputs[26][58] , 
        \negative_inputs[26][57] , \negative_inputs[26][56] , 
        \negative_inputs[26][55] , \negative_inputs[26][54] , 
        \negative_inputs[26][53] , \negative_inputs[26][52] , 
        \negative_inputs[26][51] , \negative_inputs[26][50] , 
        \negative_inputs[26][49] , \negative_inputs[26][48] , 
        \negative_inputs[26][47] , \negative_inputs[26][46] , 
        \negative_inputs[26][45] , \negative_inputs[26][44] , 
        \negative_inputs[26][43] , \negative_inputs[26][42] , 
        \negative_inputs[26][41] , \negative_inputs[26][40] , 
        \negative_inputs[26][39] , \negative_inputs[26][38] , 
        \negative_inputs[26][37] , \negative_inputs[26][36] , 
        \negative_inputs[26][35] , \negative_inputs[26][34] , 
        \negative_inputs[26][33] , \negative_inputs[26][32] , 
        \negative_inputs[26][31] , \negative_inputs[26][30] , 
        \negative_inputs[26][29] , \negative_inputs[26][28] , 
        \negative_inputs[26][27] , \negative_inputs[26][26] , 
        \negative_inputs[26][25] , \negative_inputs[26][24] , 
        \negative_inputs[26][23] , \negative_inputs[26][22] , 
        \negative_inputs[26][21] , \negative_inputs[26][20] , 
        \negative_inputs[26][19] , \negative_inputs[26][18] , 
        \negative_inputs[26][17] , \negative_inputs[26][16] , 
        \negative_inputs[26][15] , \negative_inputs[26][14] , 
        \negative_inputs[26][13] , \negative_inputs[26][12] , 
        \negative_inputs[26][11] , \negative_inputs[26][10] , 
        \negative_inputs[26][9] , \negative_inputs[26][8] , 
        \negative_inputs[26][7] , \negative_inputs[26][6] , 
        \negative_inputs[26][5] , \negative_inputs[26][4] , 
        \negative_inputs[26][3] , \negative_inputs[26][2] , 
        \negative_inputs[26][1] , \negative_inputs[26][0] }) );
  complement_NBIT64_5 complement_A_signal_27 ( .A({n656, n654, n674, n647, 
        n641, n645, n626, n623, n617, n614, n611, n609, n604, n600, n596, n593, 
        n586, n580, n574, n571, n565, n561, n555, n553, n549, n545, n540, n538, 
        n535, n531, n491, n501, n505, n495, n503, n514, n498, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[27][63] , \negative_inputs[27][62] , 
        \negative_inputs[27][61] , \negative_inputs[27][60] , 
        \negative_inputs[27][59] , \negative_inputs[27][58] , 
        \negative_inputs[27][57] , \negative_inputs[27][56] , 
        \negative_inputs[27][55] , \negative_inputs[27][54] , 
        \negative_inputs[27][53] , \negative_inputs[27][52] , 
        \negative_inputs[27][51] , \negative_inputs[27][50] , 
        \negative_inputs[27][49] , \negative_inputs[27][48] , 
        \negative_inputs[27][47] , \negative_inputs[27][46] , 
        \negative_inputs[27][45] , \negative_inputs[27][44] , 
        \negative_inputs[27][43] , \negative_inputs[27][42] , 
        \negative_inputs[27][41] , \negative_inputs[27][40] , 
        \negative_inputs[27][39] , \negative_inputs[27][38] , 
        \negative_inputs[27][37] , \negative_inputs[27][36] , 
        \negative_inputs[27][35] , \negative_inputs[27][34] , 
        \negative_inputs[27][33] , \negative_inputs[27][32] , 
        \negative_inputs[27][31] , \negative_inputs[27][30] , 
        \negative_inputs[27][29] , \negative_inputs[27][28] , 
        \negative_inputs[27][27] , \negative_inputs[27][26] , 
        \negative_inputs[27][25] , \negative_inputs[27][24] , 
        \negative_inputs[27][23] , \negative_inputs[27][22] , 
        \negative_inputs[27][21] , \negative_inputs[27][20] , 
        \negative_inputs[27][19] , \negative_inputs[27][18] , 
        \negative_inputs[27][17] , \negative_inputs[27][16] , 
        \negative_inputs[27][15] , \negative_inputs[27][14] , 
        \negative_inputs[27][13] , \negative_inputs[27][12] , 
        \negative_inputs[27][11] , \negative_inputs[27][10] , 
        \negative_inputs[27][9] , \negative_inputs[27][8] , 
        \negative_inputs[27][7] , \negative_inputs[27][6] , 
        \negative_inputs[27][5] , \negative_inputs[27][4] , 
        \negative_inputs[27][3] , \negative_inputs[27][2] , 
        \negative_inputs[27][1] , \negative_inputs[27][0] }) );
  complement_NBIT64_4 complement_A_signal_28 ( .A({n656, n654, n674, n647, 
        n641, n627, n623, n618, n614, n611, n608, n605, n599, n596, n592, n587, 
        n579, n574, n570, n566, n561, n556, n552, n550, n545, n540, n538, n535, 
        n531, n491, n490, n496, n500, n504, n513, n507, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[28][63] , \negative_inputs[28][62] , 
        \negative_inputs[28][61] , \negative_inputs[28][60] , 
        \negative_inputs[28][59] , \negative_inputs[28][58] , 
        \negative_inputs[28][57] , \negative_inputs[28][56] , 
        \negative_inputs[28][55] , \negative_inputs[28][54] , 
        \negative_inputs[28][53] , \negative_inputs[28][52] , 
        \negative_inputs[28][51] , \negative_inputs[28][50] , 
        \negative_inputs[28][49] , \negative_inputs[28][48] , 
        \negative_inputs[28][47] , \negative_inputs[28][46] , 
        \negative_inputs[28][45] , \negative_inputs[28][44] , 
        \negative_inputs[28][43] , \negative_inputs[28][42] , 
        \negative_inputs[28][41] , \negative_inputs[28][40] , 
        \negative_inputs[28][39] , \negative_inputs[28][38] , 
        \negative_inputs[28][37] , \negative_inputs[28][36] , 
        \negative_inputs[28][35] , \negative_inputs[28][34] , 
        \negative_inputs[28][33] , \negative_inputs[28][32] , 
        \negative_inputs[28][31] , \negative_inputs[28][30] , 
        \negative_inputs[28][29] , \negative_inputs[28][28] , 
        \negative_inputs[28][27] , \negative_inputs[28][26] , 
        \negative_inputs[28][25] , \negative_inputs[28][24] , 
        \negative_inputs[28][23] , \negative_inputs[28][22] , 
        \negative_inputs[28][21] , \negative_inputs[28][20] , 
        \negative_inputs[28][19] , \negative_inputs[28][18] , 
        \negative_inputs[28][17] , \negative_inputs[28][16] , 
        \negative_inputs[28][15] , \negative_inputs[28][14] , 
        \negative_inputs[28][13] , \negative_inputs[28][12] , 
        \negative_inputs[28][11] , \negative_inputs[28][10] , 
        \negative_inputs[28][9] , \negative_inputs[28][8] , 
        \negative_inputs[28][7] , \negative_inputs[28][6] , 
        \negative_inputs[28][5] , \negative_inputs[28][4] , 
        \negative_inputs[28][3] , \negative_inputs[28][2] , 
        \negative_inputs[28][1] , \negative_inputs[28][0] }) );
  complement_NBIT64_3 complement_A_signal_29 ( .A({n656, n654, n674, n647, 
        n626, n623, n617, n615, n611, n608, n604, n600, n596, n593, n586, n581, 
        n574, n571, n565, n562, n555, n553, n549, n545, n540, n538, n534, n532, 
        n491, n501, n506, n494, n504, n514, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[29][63] , \negative_inputs[29][62] , 
        \negative_inputs[29][61] , \negative_inputs[29][60] , 
        \negative_inputs[29][59] , \negative_inputs[29][58] , 
        \negative_inputs[29][57] , \negative_inputs[29][56] , 
        \negative_inputs[29][55] , \negative_inputs[29][54] , 
        \negative_inputs[29][53] , \negative_inputs[29][52] , 
        \negative_inputs[29][51] , \negative_inputs[29][50] , 
        \negative_inputs[29][49] , \negative_inputs[29][48] , 
        \negative_inputs[29][47] , \negative_inputs[29][46] , 
        \negative_inputs[29][45] , \negative_inputs[29][44] , 
        \negative_inputs[29][43] , \negative_inputs[29][42] , 
        \negative_inputs[29][41] , \negative_inputs[29][40] , 
        \negative_inputs[29][39] , \negative_inputs[29][38] , 
        \negative_inputs[29][37] , \negative_inputs[29][36] , 
        \negative_inputs[29][35] , \negative_inputs[29][34] , 
        \negative_inputs[29][33] , \negative_inputs[29][32] , 
        \negative_inputs[29][31] , \negative_inputs[29][30] , 
        \negative_inputs[29][29] , \negative_inputs[29][28] , 
        \negative_inputs[29][27] , \negative_inputs[29][26] , 
        \negative_inputs[29][25] , \negative_inputs[29][24] , 
        \negative_inputs[29][23] , \negative_inputs[29][22] , 
        \negative_inputs[29][21] , \negative_inputs[29][20] , 
        \negative_inputs[29][19] , \negative_inputs[29][18] , 
        \negative_inputs[29][17] , \negative_inputs[29][16] , 
        \negative_inputs[29][15] , \negative_inputs[29][14] , 
        \negative_inputs[29][13] , \negative_inputs[29][12] , 
        \negative_inputs[29][11] , \negative_inputs[29][10] , 
        \negative_inputs[29][9] , \negative_inputs[29][8] , 
        \negative_inputs[29][7] , \negative_inputs[29][6] , 
        \negative_inputs[29][5] , \negative_inputs[29][4] , 
        \negative_inputs[29][3] , \negative_inputs[29][2] , 
        \negative_inputs[29][1] , \negative_inputs[29][0] }) );
  complement_NBIT64_2 complement_A_signal_30 ( .A({n656, n653, n674, n627, 
        n622, n618, n614, n612, n608, n605, n599, n597, n592, n587, n579, n575, 
        n570, n565, n560, n556, n552, n550, n545, n541, n537, n535, n532, n530, 
        n490, n506, n499, n504, n513, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[30][63] , \negative_inputs[30][62] , 
        \negative_inputs[30][61] , \negative_inputs[30][60] , 
        \negative_inputs[30][59] , \negative_inputs[30][58] , 
        \negative_inputs[30][57] , \negative_inputs[30][56] , 
        \negative_inputs[30][55] , \negative_inputs[30][54] , 
        \negative_inputs[30][53] , \negative_inputs[30][52] , 
        \negative_inputs[30][51] , \negative_inputs[30][50] , 
        \negative_inputs[30][49] , \negative_inputs[30][48] , 
        \negative_inputs[30][47] , \negative_inputs[30][46] , 
        \negative_inputs[30][45] , \negative_inputs[30][44] , 
        \negative_inputs[30][43] , \negative_inputs[30][42] , 
        \negative_inputs[30][41] , \negative_inputs[30][40] , 
        \negative_inputs[30][39] , \negative_inputs[30][38] , 
        \negative_inputs[30][37] , \negative_inputs[30][36] , 
        \negative_inputs[30][35] , \negative_inputs[30][34] , 
        \negative_inputs[30][33] , \negative_inputs[30][32] , 
        \negative_inputs[30][31] , \negative_inputs[30][30] , 
        \negative_inputs[30][29] , \negative_inputs[30][28] , 
        \negative_inputs[30][27] , \negative_inputs[30][26] , 
        \negative_inputs[30][25] , \negative_inputs[30][24] , 
        \negative_inputs[30][23] , \negative_inputs[30][22] , 
        \negative_inputs[30][21] , \negative_inputs[30][20] , 
        \negative_inputs[30][19] , \negative_inputs[30][18] , 
        \negative_inputs[30][17] , \negative_inputs[30][16] , 
        \negative_inputs[30][15] , \negative_inputs[30][14] , 
        \negative_inputs[30][13] , \negative_inputs[30][12] , 
        \negative_inputs[30][11] , \negative_inputs[30][10] , 
        \negative_inputs[30][9] , \negative_inputs[30][8] , 
        \negative_inputs[30][7] , \negative_inputs[30][6] , 
        \negative_inputs[30][5] , \negative_inputs[30][4] , 
        \negative_inputs[30][3] , \negative_inputs[30][2] , 
        \negative_inputs[30][1] , \negative_inputs[30][0] }) );
  complement_NBIT64_1 complement_A_signal_31 ( .A({n656, n653, n628, n623, 
        n617, n615, n611, n609, n604, n600, n596, n593, n586, n580, n574, n571, 
        n565, n561, n555, n553, n549, n545, n540, n538, n535, n532, n491, n501, 
        n506, n520, n503, n514, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\negative_inputs[31][63] , \negative_inputs[31][62] , 
        \negative_inputs[31][61] , \negative_inputs[31][60] , 
        \negative_inputs[31][59] , \negative_inputs[31][58] , 
        \negative_inputs[31][57] , \negative_inputs[31][56] , 
        \negative_inputs[31][55] , \negative_inputs[31][54] , 
        \negative_inputs[31][53] , \negative_inputs[31][52] , 
        \negative_inputs[31][51] , \negative_inputs[31][50] , 
        \negative_inputs[31][49] , \negative_inputs[31][48] , 
        \negative_inputs[31][47] , \negative_inputs[31][46] , 
        \negative_inputs[31][45] , \negative_inputs[31][44] , 
        \negative_inputs[31][43] , \negative_inputs[31][42] , 
        \negative_inputs[31][41] , \negative_inputs[31][40] , 
        \negative_inputs[31][39] , \negative_inputs[31][38] , 
        \negative_inputs[31][37] , \negative_inputs[31][36] , 
        \negative_inputs[31][35] , \negative_inputs[31][34] , 
        \negative_inputs[31][33] , \negative_inputs[31][32] , 
        \negative_inputs[31][31] , \negative_inputs[31][30] , 
        \negative_inputs[31][29] , \negative_inputs[31][28] , 
        \negative_inputs[31][27] , \negative_inputs[31][26] , 
        \negative_inputs[31][25] , \negative_inputs[31][24] , 
        \negative_inputs[31][23] , \negative_inputs[31][22] , 
        \negative_inputs[31][21] , \negative_inputs[31][20] , 
        \negative_inputs[31][19] , \negative_inputs[31][18] , 
        \negative_inputs[31][17] , \negative_inputs[31][16] , 
        \negative_inputs[31][15] , \negative_inputs[31][14] , 
        \negative_inputs[31][13] , \negative_inputs[31][12] , 
        \negative_inputs[31][11] , \negative_inputs[31][10] , 
        \negative_inputs[31][9] , \negative_inputs[31][8] , 
        \negative_inputs[31][7] , \negative_inputs[31][6] , 
        \negative_inputs[31][5] , \negative_inputs[31][4] , 
        \negative_inputs[31][3] , \negative_inputs[31][2] , 
        \negative_inputs[31][1] , \negative_inputs[31][0] }) );
  booth_encoder_NBIT32 BOOTH_enc ( .A(in_2), .Y(Encoder_out) );
  MUX81_GENERIC_NBIT64_0 MUX81_N_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n657, 
        n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, 
        n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, n658, 
        n658, n658, n658, n658, n658, n658, n658, n659, n627, n624, n618, n615, 
        n612, n609, n606, n600, n597, n594, n587, n582, n575, n571, n566, n563, 
        n556, n553, n550, n547, n541, n537, n535, n532, n530, n527, n496, n521, 
        n517, n515, n507}), .C({n659, n659, n659, n659, n659, n659, n659, n659, 
        n659, n659, n659, n657, n659, n659, n659, n659, n659, n659, n659, n659, 
        n659, n659, n659, n659, n658, n659, n659, n659, n659, n659, n659, n659, 
        n627, n624, n618, n615, n612, n609, n606, n600, n597, n593, n587, n582, 
        n575, n571, n566, n563, n556, n553, n550, n547, n541, n538, n534, n532, 
        n530, n527, n496, n520, n518, n514, n507, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[0][63] , \negative_inputs[0][62] , 
        \negative_inputs[0][61] , \negative_inputs[0][60] , 
        \negative_inputs[0][59] , \negative_inputs[0][58] , 
        \negative_inputs[0][57] , \negative_inputs[0][56] , 
        \negative_inputs[0][55] , \negative_inputs[0][54] , 
        \negative_inputs[0][53] , \negative_inputs[0][52] , 
        \negative_inputs[0][51] , \negative_inputs[0][50] , 
        \negative_inputs[0][49] , \negative_inputs[0][48] , 
        \negative_inputs[0][47] , \negative_inputs[0][46] , 
        \negative_inputs[0][45] , \negative_inputs[0][44] , 
        \negative_inputs[0][43] , \negative_inputs[0][42] , 
        \negative_inputs[0][41] , \negative_inputs[0][40] , 
        \negative_inputs[0][39] , \negative_inputs[0][38] , 
        \negative_inputs[0][37] , \negative_inputs[0][36] , 
        \negative_inputs[0][35] , \negative_inputs[0][34] , 
        \negative_inputs[0][33] , \negative_inputs[0][32] , 
        \negative_inputs[0][31] , \negative_inputs[0][30] , 
        \negative_inputs[0][29] , \negative_inputs[0][28] , 
        \negative_inputs[0][27] , \negative_inputs[0][26] , 
        \negative_inputs[0][25] , \negative_inputs[0][24] , 
        \negative_inputs[0][23] , \negative_inputs[0][22] , 
        \negative_inputs[0][21] , \negative_inputs[0][20] , 
        \negative_inputs[0][19] , \negative_inputs[0][18] , 
        \negative_inputs[0][17] , \negative_inputs[0][16] , 
        \negative_inputs[0][15] , \negative_inputs[0][14] , 
        \negative_inputs[0][13] , \negative_inputs[0][12] , 
        \negative_inputs[0][11] , \negative_inputs[0][10] , 
        \negative_inputs[0][9] , \negative_inputs[0][8] , 
        \negative_inputs[0][7] , \negative_inputs[0][6] , 
        \negative_inputs[0][5] , \negative_inputs[0][4] , 
        \negative_inputs[0][3] , \negative_inputs[0][2] , 
        \negative_inputs[0][1] , \negative_inputs[0][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[1][63] , \negative_inputs[1][62] , 
        \negative_inputs[1][61] , \negative_inputs[1][60] , 
        \negative_inputs[1][59] , \negative_inputs[1][58] , 
        \negative_inputs[1][57] , \negative_inputs[1][56] , 
        \negative_inputs[1][55] , \negative_inputs[1][54] , 
        \negative_inputs[1][53] , \negative_inputs[1][52] , 
        \negative_inputs[1][51] , \negative_inputs[1][50] , 
        \negative_inputs[1][49] , \negative_inputs[1][48] , 
        \negative_inputs[1][47] , \negative_inputs[1][46] , 
        \negative_inputs[1][45] , \negative_inputs[1][44] , 
        \negative_inputs[1][43] , \negative_inputs[1][42] , 
        \negative_inputs[1][41] , \negative_inputs[1][40] , 
        \negative_inputs[1][39] , \negative_inputs[1][38] , 
        \negative_inputs[1][37] , \negative_inputs[1][36] , 
        \negative_inputs[1][35] , \negative_inputs[1][34] , 
        \negative_inputs[1][33] , \negative_inputs[1][32] , 
        \negative_inputs[1][31] , \negative_inputs[1][30] , 
        \negative_inputs[1][29] , \negative_inputs[1][28] , 
        \negative_inputs[1][27] , \negative_inputs[1][26] , 
        \negative_inputs[1][25] , \negative_inputs[1][24] , 
        \negative_inputs[1][23] , \negative_inputs[1][22] , 
        \negative_inputs[1][21] , \negative_inputs[1][20] , 
        \negative_inputs[1][19] , \negative_inputs[1][18] , 
        \negative_inputs[1][17] , \negative_inputs[1][16] , 
        \negative_inputs[1][15] , \negative_inputs[1][14] , 
        \negative_inputs[1][13] , \negative_inputs[1][12] , 
        \negative_inputs[1][11] , \negative_inputs[1][10] , 
        \negative_inputs[1][9] , \negative_inputs[1][8] , 
        \negative_inputs[1][7] , \negative_inputs[1][6] , 
        \negative_inputs[1][5] , \negative_inputs[1][4] , 
        \negative_inputs[1][3] , \negative_inputs[1][2] , 
        \negative_inputs[1][1] , \negative_inputs[1][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[2:0]), .Y({\ADDER_IN_from_mux[0][63] , 
        \ADDER_IN_from_mux[0][62] , \ADDER_IN_from_mux[0][61] , 
        \ADDER_IN_from_mux[0][60] , \ADDER_IN_from_mux[0][59] , 
        \ADDER_IN_from_mux[0][58] , \ADDER_IN_from_mux[0][57] , 
        \ADDER_IN_from_mux[0][56] , \ADDER_IN_from_mux[0][55] , 
        \ADDER_IN_from_mux[0][54] , \ADDER_IN_from_mux[0][53] , 
        \ADDER_IN_from_mux[0][52] , \ADDER_IN_from_mux[0][51] , 
        \ADDER_IN_from_mux[0][50] , \ADDER_IN_from_mux[0][49] , 
        \ADDER_IN_from_mux[0][48] , \ADDER_IN_from_mux[0][47] , 
        \ADDER_IN_from_mux[0][46] , \ADDER_IN_from_mux[0][45] , 
        \ADDER_IN_from_mux[0][44] , \ADDER_IN_from_mux[0][43] , 
        \ADDER_IN_from_mux[0][42] , \ADDER_IN_from_mux[0][41] , 
        \ADDER_IN_from_mux[0][40] , \ADDER_IN_from_mux[0][39] , 
        \ADDER_IN_from_mux[0][38] , \ADDER_IN_from_mux[0][37] , 
        \ADDER_IN_from_mux[0][36] , \ADDER_IN_from_mux[0][35] , 
        \ADDER_IN_from_mux[0][34] , \ADDER_IN_from_mux[0][33] , 
        \ADDER_IN_from_mux[0][32] , \ADDER_IN_from_mux[0][31] , 
        \ADDER_IN_from_mux[0][30] , \ADDER_IN_from_mux[0][29] , 
        \ADDER_IN_from_mux[0][28] , \ADDER_IN_from_mux[0][27] , 
        \ADDER_IN_from_mux[0][26] , \ADDER_IN_from_mux[0][25] , 
        \ADDER_IN_from_mux[0][24] , \ADDER_IN_from_mux[0][23] , 
        \ADDER_IN_from_mux[0][22] , \ADDER_IN_from_mux[0][21] , 
        \ADDER_IN_from_mux[0][20] , \ADDER_IN_from_mux[0][19] , 
        \ADDER_IN_from_mux[0][18] , \ADDER_IN_from_mux[0][17] , 
        \ADDER_IN_from_mux[0][16] , \ADDER_IN_from_mux[0][15] , 
        \ADDER_IN_from_mux[0][14] , \ADDER_IN_from_mux[0][13] , 
        \ADDER_IN_from_mux[0][12] , \ADDER_IN_from_mux[0][11] , 
        \ADDER_IN_from_mux[0][10] , \ADDER_IN_from_mux[0][9] , 
        \ADDER_IN_from_mux[0][8] , \ADDER_IN_from_mux[0][7] , 
        \ADDER_IN_from_mux[0][6] , \ADDER_IN_from_mux[0][5] , 
        \ADDER_IN_from_mux[0][4] , \ADDER_IN_from_mux[0][3] , 
        \ADDER_IN_from_mux[0][2] , \ADDER_IN_from_mux[0][1] , 
        \ADDER_IN_from_mux[0][0] }) );
  MUX81_GENERIC_NBIT64_15 MUX81_N_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n670, 
        n670, n670, n670, n670, n671, n671, n671, n671, n671, n671, n671, n671, 
        n671, n671, n671, n671, n671, n671, n671, n671, n671, n671, n671, n671, 
        n671, n671, n672, n672, n672, n672, n628, n625, n619, n616, n613, n610, 
        n606, n601, n598, n594, n588, n582, n576, n572, n567, n563, n557, n554, 
        n551, n547, n542, n537, n535, n532, n530, n527, n506, n521, n517, n515, 
        n507, 1'b0, 1'b0}), .C({n657, n657, n658, n657, n657, n657, n657, n658, 
        n657, n657, n657, n657, n657, n657, n657, n657, n658, n664, n663, n663, 
        n663, n663, n663, n663, n663, n663, n663, n663, n663, n663, n627, n624, 
        n618, n615, n612, n609, n606, n600, n597, n594, n587, n582, n575, n571, 
        n566, n563, n556, n553, n550, n547, n541, n537, n535, n532, n530, n527, 
        n496, n495, n517, n515, n507, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[2][63] , \negative_inputs[2][62] , 
        \negative_inputs[2][61] , \negative_inputs[2][60] , 
        \negative_inputs[2][59] , \negative_inputs[2][58] , 
        \negative_inputs[2][57] , \negative_inputs[2][56] , 
        \negative_inputs[2][55] , \negative_inputs[2][54] , 
        \negative_inputs[2][53] , \negative_inputs[2][52] , 
        \negative_inputs[2][51] , \negative_inputs[2][50] , 
        \negative_inputs[2][49] , \negative_inputs[2][48] , 
        \negative_inputs[2][47] , \negative_inputs[2][46] , 
        \negative_inputs[2][45] , \negative_inputs[2][44] , 
        \negative_inputs[2][43] , \negative_inputs[2][42] , 
        \negative_inputs[2][41] , \negative_inputs[2][40] , 
        \negative_inputs[2][39] , \negative_inputs[2][38] , 
        \negative_inputs[2][37] , \negative_inputs[2][36] , 
        \negative_inputs[2][35] , \negative_inputs[2][34] , 
        \negative_inputs[2][33] , \negative_inputs[2][32] , 
        \negative_inputs[2][31] , \negative_inputs[2][30] , 
        \negative_inputs[2][29] , \negative_inputs[2][28] , 
        \negative_inputs[2][27] , \negative_inputs[2][26] , 
        \negative_inputs[2][25] , \negative_inputs[2][24] , 
        \negative_inputs[2][23] , \negative_inputs[2][22] , 
        \negative_inputs[2][21] , \negative_inputs[2][20] , 
        \negative_inputs[2][19] , \negative_inputs[2][18] , 
        \negative_inputs[2][17] , \negative_inputs[2][16] , 
        \negative_inputs[2][15] , \negative_inputs[2][14] , 
        \negative_inputs[2][13] , \negative_inputs[2][12] , 
        \negative_inputs[2][11] , \negative_inputs[2][10] , 
        \negative_inputs[2][9] , \negative_inputs[2][8] , 
        \negative_inputs[2][7] , \negative_inputs[2][6] , 
        \negative_inputs[2][5] , \negative_inputs[2][4] , 
        \negative_inputs[2][3] , \negative_inputs[2][2] , 
        \negative_inputs[2][1] , \negative_inputs[2][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[3][63] , \negative_inputs[3][62] , 
        \negative_inputs[3][61] , \negative_inputs[3][60] , 
        \negative_inputs[3][59] , \negative_inputs[3][58] , 
        \negative_inputs[3][57] , \negative_inputs[3][56] , 
        \negative_inputs[3][55] , \negative_inputs[3][54] , 
        \negative_inputs[3][53] , \negative_inputs[3][52] , 
        \negative_inputs[3][51] , \negative_inputs[3][50] , 
        \negative_inputs[3][49] , \negative_inputs[3][48] , 
        \negative_inputs[3][47] , \negative_inputs[3][46] , 
        \negative_inputs[3][45] , \negative_inputs[3][44] , 
        \negative_inputs[3][43] , \negative_inputs[3][42] , 
        \negative_inputs[3][41] , \negative_inputs[3][40] , 
        \negative_inputs[3][39] , \negative_inputs[3][38] , 
        \negative_inputs[3][37] , \negative_inputs[3][36] , 
        \negative_inputs[3][35] , \negative_inputs[3][34] , 
        \negative_inputs[3][33] , \negative_inputs[3][32] , 
        \negative_inputs[3][31] , \negative_inputs[3][30] , 
        \negative_inputs[3][29] , \negative_inputs[3][28] , 
        \negative_inputs[3][27] , \negative_inputs[3][26] , 
        \negative_inputs[3][25] , \negative_inputs[3][24] , 
        \negative_inputs[3][23] , \negative_inputs[3][22] , 
        \negative_inputs[3][21] , \negative_inputs[3][20] , 
        \negative_inputs[3][19] , \negative_inputs[3][18] , 
        \negative_inputs[3][17] , \negative_inputs[3][16] , 
        \negative_inputs[3][15] , \negative_inputs[3][14] , 
        \negative_inputs[3][13] , \negative_inputs[3][12] , 
        \negative_inputs[3][11] , \negative_inputs[3][10] , 
        \negative_inputs[3][9] , \negative_inputs[3][8] , 
        \negative_inputs[3][7] , \negative_inputs[3][6] , 
        \negative_inputs[3][5] , \negative_inputs[3][4] , 
        \negative_inputs[3][3] , \negative_inputs[3][2] , 
        \negative_inputs[3][1] , \negative_inputs[3][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[5:3]), .Y({\ADDER_IN_from_mux[1][63] , 
        \ADDER_IN_from_mux[1][62] , \ADDER_IN_from_mux[1][61] , 
        \ADDER_IN_from_mux[1][60] , \ADDER_IN_from_mux[1][59] , 
        \ADDER_IN_from_mux[1][58] , \ADDER_IN_from_mux[1][57] , 
        \ADDER_IN_from_mux[1][56] , \ADDER_IN_from_mux[1][55] , 
        \ADDER_IN_from_mux[1][54] , \ADDER_IN_from_mux[1][53] , 
        \ADDER_IN_from_mux[1][52] , \ADDER_IN_from_mux[1][51] , 
        \ADDER_IN_from_mux[1][50] , \ADDER_IN_from_mux[1][49] , 
        \ADDER_IN_from_mux[1][48] , \ADDER_IN_from_mux[1][47] , 
        \ADDER_IN_from_mux[1][46] , \ADDER_IN_from_mux[1][45] , 
        \ADDER_IN_from_mux[1][44] , \ADDER_IN_from_mux[1][43] , 
        \ADDER_IN_from_mux[1][42] , \ADDER_IN_from_mux[1][41] , 
        \ADDER_IN_from_mux[1][40] , \ADDER_IN_from_mux[1][39] , 
        \ADDER_IN_from_mux[1][38] , \ADDER_IN_from_mux[1][37] , 
        \ADDER_IN_from_mux[1][36] , \ADDER_IN_from_mux[1][35] , 
        \ADDER_IN_from_mux[1][34] , \ADDER_IN_from_mux[1][33] , 
        \ADDER_IN_from_mux[1][32] , \ADDER_IN_from_mux[1][31] , 
        \ADDER_IN_from_mux[1][30] , \ADDER_IN_from_mux[1][29] , 
        \ADDER_IN_from_mux[1][28] , \ADDER_IN_from_mux[1][27] , 
        \ADDER_IN_from_mux[1][26] , \ADDER_IN_from_mux[1][25] , 
        \ADDER_IN_from_mux[1][24] , \ADDER_IN_from_mux[1][23] , 
        \ADDER_IN_from_mux[1][22] , \ADDER_IN_from_mux[1][21] , 
        \ADDER_IN_from_mux[1][20] , \ADDER_IN_from_mux[1][19] , 
        \ADDER_IN_from_mux[1][18] , \ADDER_IN_from_mux[1][17] , 
        \ADDER_IN_from_mux[1][16] , \ADDER_IN_from_mux[1][15] , 
        \ADDER_IN_from_mux[1][14] , \ADDER_IN_from_mux[1][13] , 
        \ADDER_IN_from_mux[1][12] , \ADDER_IN_from_mux[1][11] , 
        \ADDER_IN_from_mux[1][10] , \ADDER_IN_from_mux[1][9] , 
        \ADDER_IN_from_mux[1][8] , \ADDER_IN_from_mux[1][7] , 
        \ADDER_IN_from_mux[1][6] , \ADDER_IN_from_mux[1][5] , 
        \ADDER_IN_from_mux[1][4] , \ADDER_IN_from_mux[1][3] , 
        \ADDER_IN_from_mux[1][2] , \ADDER_IN_from_mux[1][1] , 
        \ADDER_IN_from_mux[1][0] }) );
  MUX81_GENERIC_NBIT64_14 MUX81_N_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n663, 
        n663, n663, n663, n663, n663, n663, n663, n663, n663, n663, n663, n663, 
        n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, 
        n664, n664, n664, n664, n627, n624, n618, n615, n612, n609, n606, n600, 
        n597, n594, n587, n582, n575, n572, n566, n563, n556, n553, n550, n547, 
        n541, n538, n534, n532, n529, n527, n496, n521, n517, n515, n507, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n672, n672, n672, n672, n672, n672, n672, n672, 
        n673, n673, n673, n673, n673, n673, n673, n673, n673, n673, n672, n672, 
        n672, n672, n672, n672, n672, n672, n672, n672, n628, n624, n619, n616, 
        n613, n610, n606, n601, n598, n594, n588, n583, n576, n572, n567, n564, 
        n557, n554, n551, n547, n542, n537, n535, n531, n529, n527, n506, n521, 
        n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[4][63] , \negative_inputs[4][62] , 
        \negative_inputs[4][61] , \negative_inputs[4][60] , 
        \negative_inputs[4][59] , \negative_inputs[4][58] , 
        \negative_inputs[4][57] , \negative_inputs[4][56] , 
        \negative_inputs[4][55] , \negative_inputs[4][54] , 
        \negative_inputs[4][53] , \negative_inputs[4][52] , 
        \negative_inputs[4][51] , \negative_inputs[4][50] , 
        \negative_inputs[4][49] , \negative_inputs[4][48] , 
        \negative_inputs[4][47] , \negative_inputs[4][46] , 
        \negative_inputs[4][45] , \negative_inputs[4][44] , 
        \negative_inputs[4][43] , \negative_inputs[4][42] , 
        \negative_inputs[4][41] , \negative_inputs[4][40] , 
        \negative_inputs[4][39] , \negative_inputs[4][38] , 
        \negative_inputs[4][37] , \negative_inputs[4][36] , 
        \negative_inputs[4][35] , \negative_inputs[4][34] , 
        \negative_inputs[4][33] , \negative_inputs[4][32] , 
        \negative_inputs[4][31] , \negative_inputs[4][30] , 
        \negative_inputs[4][29] , \negative_inputs[4][28] , 
        \negative_inputs[4][27] , \negative_inputs[4][26] , 
        \negative_inputs[4][25] , \negative_inputs[4][24] , 
        \negative_inputs[4][23] , \negative_inputs[4][22] , 
        \negative_inputs[4][21] , \negative_inputs[4][20] , 
        \negative_inputs[4][19] , \negative_inputs[4][18] , 
        \negative_inputs[4][17] , \negative_inputs[4][16] , 
        \negative_inputs[4][15] , \negative_inputs[4][14] , 
        \negative_inputs[4][13] , \negative_inputs[4][12] , 
        \negative_inputs[4][11] , \negative_inputs[4][10] , 
        \negative_inputs[4][9] , \negative_inputs[4][8] , 
        \negative_inputs[4][7] , \negative_inputs[4][6] , 
        \negative_inputs[4][5] , \negative_inputs[4][4] , 
        \negative_inputs[4][3] , \negative_inputs[4][2] , 
        \negative_inputs[4][1] , \negative_inputs[4][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[5][63] , \negative_inputs[5][62] , 
        \negative_inputs[5][61] , \negative_inputs[5][60] , 
        \negative_inputs[5][59] , \negative_inputs[5][58] , 
        \negative_inputs[5][57] , \negative_inputs[5][56] , 
        \negative_inputs[5][55] , \negative_inputs[5][54] , 
        \negative_inputs[5][53] , \negative_inputs[5][52] , 
        \negative_inputs[5][51] , \negative_inputs[5][50] , 
        \negative_inputs[5][49] , \negative_inputs[5][48] , 
        \negative_inputs[5][47] , \negative_inputs[5][46] , 
        \negative_inputs[5][45] , \negative_inputs[5][44] , 
        \negative_inputs[5][43] , \negative_inputs[5][42] , 
        \negative_inputs[5][41] , \negative_inputs[5][40] , 
        \negative_inputs[5][39] , \negative_inputs[5][38] , 
        \negative_inputs[5][37] , \negative_inputs[5][36] , 
        \negative_inputs[5][35] , \negative_inputs[5][34] , 
        \negative_inputs[5][33] , \negative_inputs[5][32] , 
        \negative_inputs[5][31] , \negative_inputs[5][30] , 
        \negative_inputs[5][29] , \negative_inputs[5][28] , 
        \negative_inputs[5][27] , \negative_inputs[5][26] , 
        \negative_inputs[5][25] , \negative_inputs[5][24] , 
        \negative_inputs[5][23] , \negative_inputs[5][22] , 
        \negative_inputs[5][21] , \negative_inputs[5][20] , 
        \negative_inputs[5][19] , \negative_inputs[5][18] , 
        \negative_inputs[5][17] , \negative_inputs[5][16] , 
        \negative_inputs[5][15] , \negative_inputs[5][14] , 
        \negative_inputs[5][13] , \negative_inputs[5][12] , 
        \negative_inputs[5][11] , \negative_inputs[5][10] , 
        \negative_inputs[5][9] , \negative_inputs[5][8] , 
        \negative_inputs[5][7] , \negative_inputs[5][6] , 
        \negative_inputs[5][5] , \negative_inputs[5][4] , 
        \negative_inputs[5][3] , \negative_inputs[5][2] , 
        \negative_inputs[5][1] , \negative_inputs[5][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[8:6]), .Y({\ADDER_IN_from_mux[2][63] , 
        \ADDER_IN_from_mux[2][62] , \ADDER_IN_from_mux[2][61] , 
        \ADDER_IN_from_mux[2][60] , \ADDER_IN_from_mux[2][59] , 
        \ADDER_IN_from_mux[2][58] , \ADDER_IN_from_mux[2][57] , 
        \ADDER_IN_from_mux[2][56] , \ADDER_IN_from_mux[2][55] , 
        \ADDER_IN_from_mux[2][54] , \ADDER_IN_from_mux[2][53] , 
        \ADDER_IN_from_mux[2][52] , \ADDER_IN_from_mux[2][51] , 
        \ADDER_IN_from_mux[2][50] , \ADDER_IN_from_mux[2][49] , 
        \ADDER_IN_from_mux[2][48] , \ADDER_IN_from_mux[2][47] , 
        \ADDER_IN_from_mux[2][46] , \ADDER_IN_from_mux[2][45] , 
        \ADDER_IN_from_mux[2][44] , \ADDER_IN_from_mux[2][43] , 
        \ADDER_IN_from_mux[2][42] , \ADDER_IN_from_mux[2][41] , 
        \ADDER_IN_from_mux[2][40] , \ADDER_IN_from_mux[2][39] , 
        \ADDER_IN_from_mux[2][38] , \ADDER_IN_from_mux[2][37] , 
        \ADDER_IN_from_mux[2][36] , \ADDER_IN_from_mux[2][35] , 
        \ADDER_IN_from_mux[2][34] , \ADDER_IN_from_mux[2][33] , 
        \ADDER_IN_from_mux[2][32] , \ADDER_IN_from_mux[2][31] , 
        \ADDER_IN_from_mux[2][30] , \ADDER_IN_from_mux[2][29] , 
        \ADDER_IN_from_mux[2][28] , \ADDER_IN_from_mux[2][27] , 
        \ADDER_IN_from_mux[2][26] , \ADDER_IN_from_mux[2][25] , 
        \ADDER_IN_from_mux[2][24] , \ADDER_IN_from_mux[2][23] , 
        \ADDER_IN_from_mux[2][22] , \ADDER_IN_from_mux[2][21] , 
        \ADDER_IN_from_mux[2][20] , \ADDER_IN_from_mux[2][19] , 
        \ADDER_IN_from_mux[2][18] , \ADDER_IN_from_mux[2][17] , 
        \ADDER_IN_from_mux[2][16] , \ADDER_IN_from_mux[2][15] , 
        \ADDER_IN_from_mux[2][14] , \ADDER_IN_from_mux[2][13] , 
        \ADDER_IN_from_mux[2][12] , \ADDER_IN_from_mux[2][11] , 
        \ADDER_IN_from_mux[2][10] , \ADDER_IN_from_mux[2][9] , 
        \ADDER_IN_from_mux[2][8] , \ADDER_IN_from_mux[2][7] , 
        \ADDER_IN_from_mux[2][6] , \ADDER_IN_from_mux[2][5] , 
        \ADDER_IN_from_mux[2][4] , \ADDER_IN_from_mux[2][3] , 
        \ADDER_IN_from_mux[2][2] , \ADDER_IN_from_mux[2][1] , 
        \ADDER_IN_from_mux[2][0] }) );
  MUX81_GENERIC_NBIT64_13 MUX81_N_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n664, 
        n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, n664, 
        n664, n664, n664, n664, n664, n665, n665, n665, n665, n665, n665, n665, 
        n665, n665, n627, n624, n618, n615, n612, n609, n606, n600, n597, n594, 
        n588, n582, n575, n572, n566, n563, n556, n553, n550, n547, n541, n538, 
        n534, n532, n491, n527, n496, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n672, n672, n672, n672, n672, n672, n672, n672, 
        n666, n666, n666, n666, n666, n667, n667, n667, n667, n667, n667, n667, 
        n667, n667, n667, n667, n667, n667, n628, n624, n619, n616, n613, n610, 
        n606, n601, n598, n594, n588, n583, n576, n572, n567, n564, n557, n554, 
        n551, n547, n542, n538, n535, n532, n491, n527, n506, n521, n517, n515, 
        n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[6][63] , \negative_inputs[6][62] , 
        \negative_inputs[6][61] , \negative_inputs[6][60] , 
        \negative_inputs[6][59] , \negative_inputs[6][58] , 
        \negative_inputs[6][57] , \negative_inputs[6][56] , 
        \negative_inputs[6][55] , \negative_inputs[6][54] , 
        \negative_inputs[6][53] , \negative_inputs[6][52] , 
        \negative_inputs[6][51] , \negative_inputs[6][50] , 
        \negative_inputs[6][49] , \negative_inputs[6][48] , 
        \negative_inputs[6][47] , \negative_inputs[6][46] , 
        \negative_inputs[6][45] , \negative_inputs[6][44] , 
        \negative_inputs[6][43] , \negative_inputs[6][42] , 
        \negative_inputs[6][41] , \negative_inputs[6][40] , 
        \negative_inputs[6][39] , \negative_inputs[6][38] , 
        \negative_inputs[6][37] , \negative_inputs[6][36] , 
        \negative_inputs[6][35] , \negative_inputs[6][34] , 
        \negative_inputs[6][33] , \negative_inputs[6][32] , 
        \negative_inputs[6][31] , \negative_inputs[6][30] , 
        \negative_inputs[6][29] , \negative_inputs[6][28] , 
        \negative_inputs[6][27] , \negative_inputs[6][26] , 
        \negative_inputs[6][25] , \negative_inputs[6][24] , 
        \negative_inputs[6][23] , \negative_inputs[6][22] , 
        \negative_inputs[6][21] , \negative_inputs[6][20] , 
        \negative_inputs[6][19] , \negative_inputs[6][18] , 
        \negative_inputs[6][17] , \negative_inputs[6][16] , 
        \negative_inputs[6][15] , \negative_inputs[6][14] , 
        \negative_inputs[6][13] , \negative_inputs[6][12] , 
        \negative_inputs[6][11] , \negative_inputs[6][10] , 
        \negative_inputs[6][9] , \negative_inputs[6][8] , 
        \negative_inputs[6][7] , \negative_inputs[6][6] , 
        \negative_inputs[6][5] , \negative_inputs[6][4] , 
        \negative_inputs[6][3] , \negative_inputs[6][2] , 
        \negative_inputs[6][1] , \negative_inputs[6][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[7][63] , \negative_inputs[7][62] , 
        \negative_inputs[7][61] , \negative_inputs[7][60] , 
        \negative_inputs[7][59] , \negative_inputs[7][58] , 
        \negative_inputs[7][57] , \negative_inputs[7][56] , 
        \negative_inputs[7][55] , \negative_inputs[7][54] , 
        \negative_inputs[7][53] , \negative_inputs[7][52] , 
        \negative_inputs[7][51] , \negative_inputs[7][50] , 
        \negative_inputs[7][49] , \negative_inputs[7][48] , 
        \negative_inputs[7][47] , \negative_inputs[7][46] , 
        \negative_inputs[7][45] , \negative_inputs[7][44] , 
        \negative_inputs[7][43] , \negative_inputs[7][42] , 
        \negative_inputs[7][41] , \negative_inputs[7][40] , 
        \negative_inputs[7][39] , \negative_inputs[7][38] , 
        \negative_inputs[7][37] , \negative_inputs[7][36] , 
        \negative_inputs[7][35] , \negative_inputs[7][34] , 
        \negative_inputs[7][33] , \negative_inputs[7][32] , 
        \negative_inputs[7][31] , \negative_inputs[7][30] , 
        \negative_inputs[7][29] , \negative_inputs[7][28] , 
        \negative_inputs[7][27] , \negative_inputs[7][26] , 
        \negative_inputs[7][25] , \negative_inputs[7][24] , 
        \negative_inputs[7][23] , \negative_inputs[7][22] , 
        \negative_inputs[7][21] , \negative_inputs[7][20] , 
        \negative_inputs[7][19] , \negative_inputs[7][18] , 
        \negative_inputs[7][17] , \negative_inputs[7][16] , 
        \negative_inputs[7][15] , \negative_inputs[7][14] , 
        \negative_inputs[7][13] , \negative_inputs[7][12] , 
        \negative_inputs[7][11] , \negative_inputs[7][10] , 
        \negative_inputs[7][9] , \negative_inputs[7][8] , 
        \negative_inputs[7][7] , \negative_inputs[7][6] , 
        \negative_inputs[7][5] , \negative_inputs[7][4] , 
        \negative_inputs[7][3] , \negative_inputs[7][2] , 
        \negative_inputs[7][1] , \negative_inputs[7][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[11:9]), .Y({\ADDER_IN_from_mux[3][63] , 
        \ADDER_IN_from_mux[3][62] , \ADDER_IN_from_mux[3][61] , 
        \ADDER_IN_from_mux[3][60] , \ADDER_IN_from_mux[3][59] , 
        \ADDER_IN_from_mux[3][58] , \ADDER_IN_from_mux[3][57] , 
        \ADDER_IN_from_mux[3][56] , \ADDER_IN_from_mux[3][55] , 
        \ADDER_IN_from_mux[3][54] , \ADDER_IN_from_mux[3][53] , 
        \ADDER_IN_from_mux[3][52] , \ADDER_IN_from_mux[3][51] , 
        \ADDER_IN_from_mux[3][50] , \ADDER_IN_from_mux[3][49] , 
        \ADDER_IN_from_mux[3][48] , \ADDER_IN_from_mux[3][47] , 
        \ADDER_IN_from_mux[3][46] , \ADDER_IN_from_mux[3][45] , 
        \ADDER_IN_from_mux[3][44] , \ADDER_IN_from_mux[3][43] , 
        \ADDER_IN_from_mux[3][42] , \ADDER_IN_from_mux[3][41] , 
        \ADDER_IN_from_mux[3][40] , \ADDER_IN_from_mux[3][39] , 
        \ADDER_IN_from_mux[3][38] , \ADDER_IN_from_mux[3][37] , 
        \ADDER_IN_from_mux[3][36] , \ADDER_IN_from_mux[3][35] , 
        \ADDER_IN_from_mux[3][34] , \ADDER_IN_from_mux[3][33] , 
        \ADDER_IN_from_mux[3][32] , \ADDER_IN_from_mux[3][31] , 
        \ADDER_IN_from_mux[3][30] , \ADDER_IN_from_mux[3][29] , 
        \ADDER_IN_from_mux[3][28] , \ADDER_IN_from_mux[3][27] , 
        \ADDER_IN_from_mux[3][26] , \ADDER_IN_from_mux[3][25] , 
        \ADDER_IN_from_mux[3][24] , \ADDER_IN_from_mux[3][23] , 
        \ADDER_IN_from_mux[3][22] , \ADDER_IN_from_mux[3][21] , 
        \ADDER_IN_from_mux[3][20] , \ADDER_IN_from_mux[3][19] , 
        \ADDER_IN_from_mux[3][18] , \ADDER_IN_from_mux[3][17] , 
        \ADDER_IN_from_mux[3][16] , \ADDER_IN_from_mux[3][15] , 
        \ADDER_IN_from_mux[3][14] , \ADDER_IN_from_mux[3][13] , 
        \ADDER_IN_from_mux[3][12] , \ADDER_IN_from_mux[3][11] , 
        \ADDER_IN_from_mux[3][10] , \ADDER_IN_from_mux[3][9] , 
        \ADDER_IN_from_mux[3][8] , \ADDER_IN_from_mux[3][7] , 
        \ADDER_IN_from_mux[3][6] , \ADDER_IN_from_mux[3][5] , 
        \ADDER_IN_from_mux[3][4] , \ADDER_IN_from_mux[3][3] , 
        \ADDER_IN_from_mux[3][2] , \ADDER_IN_from_mux[3][1] , 
        \ADDER_IN_from_mux[3][0] }) );
  MUX81_GENERIC_NBIT64_12 MUX81_N_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n665, 
        n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, 
        n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, n665, 
        n627, n624, n618, n616, n612, n609, n606, n601, n597, n594, n588, n582, 
        n575, n572, n566, n563, n556, n553, n550, n547, n541, n538, n535, n532, 
        n491, n527, n496, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n667, n667, n667, n667, n667, n667, n667, n667, 
        n667, n667, n667, n667, n667, n668, n668, n668, n668, n668, n668, n668, 
        n668, n668, n668, n668, n628, n624, n619, n616, n613, n610, n606, n601, 
        n598, n594, n588, n583, n576, n572, n567, n564, n557, n554, n551, n547, 
        n542, n538, n535, n532, n491, n527, n506, n521, n517, n515, n493, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[8][63] , \negative_inputs[8][62] , 
        \negative_inputs[8][61] , \negative_inputs[8][60] , 
        \negative_inputs[8][59] , \negative_inputs[8][58] , 
        \negative_inputs[8][57] , \negative_inputs[8][56] , 
        \negative_inputs[8][55] , \negative_inputs[8][54] , 
        \negative_inputs[8][53] , \negative_inputs[8][52] , 
        \negative_inputs[8][51] , \negative_inputs[8][50] , 
        \negative_inputs[8][49] , \negative_inputs[8][48] , 
        \negative_inputs[8][47] , \negative_inputs[8][46] , 
        \negative_inputs[8][45] , \negative_inputs[8][44] , 
        \negative_inputs[8][43] , \negative_inputs[8][42] , 
        \negative_inputs[8][41] , \negative_inputs[8][40] , 
        \negative_inputs[8][39] , \negative_inputs[8][38] , 
        \negative_inputs[8][37] , \negative_inputs[8][36] , 
        \negative_inputs[8][35] , \negative_inputs[8][34] , 
        \negative_inputs[8][33] , \negative_inputs[8][32] , 
        \negative_inputs[8][31] , \negative_inputs[8][30] , 
        \negative_inputs[8][29] , \negative_inputs[8][28] , 
        \negative_inputs[8][27] , \negative_inputs[8][26] , 
        \negative_inputs[8][25] , \negative_inputs[8][24] , 
        \negative_inputs[8][23] , \negative_inputs[8][22] , 
        \negative_inputs[8][21] , \negative_inputs[8][20] , 
        \negative_inputs[8][19] , \negative_inputs[8][18] , 
        \negative_inputs[8][17] , \negative_inputs[8][16] , 
        \negative_inputs[8][15] , \negative_inputs[8][14] , 
        \negative_inputs[8][13] , \negative_inputs[8][12] , 
        \negative_inputs[8][11] , \negative_inputs[8][10] , 
        \negative_inputs[8][9] , \negative_inputs[8][8] , 
        \negative_inputs[8][7] , \negative_inputs[8][6] , 
        \negative_inputs[8][5] , \negative_inputs[8][4] , 
        \negative_inputs[8][3] , \negative_inputs[8][2] , 
        \negative_inputs[8][1] , \negative_inputs[8][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[9][63] , \negative_inputs[9][62] , 
        \negative_inputs[9][61] , \negative_inputs[9][60] , 
        \negative_inputs[9][59] , \negative_inputs[9][58] , 
        \negative_inputs[9][57] , \negative_inputs[9][56] , 
        \negative_inputs[9][55] , \negative_inputs[9][54] , 
        \negative_inputs[9][53] , \negative_inputs[9][52] , 
        \negative_inputs[9][51] , \negative_inputs[9][50] , 
        \negative_inputs[9][49] , \negative_inputs[9][48] , 
        \negative_inputs[9][47] , \negative_inputs[9][46] , 
        \negative_inputs[9][45] , \negative_inputs[9][44] , 
        \negative_inputs[9][43] , \negative_inputs[9][42] , 
        \negative_inputs[9][41] , \negative_inputs[9][40] , 
        \negative_inputs[9][39] , \negative_inputs[9][38] , 
        \negative_inputs[9][37] , \negative_inputs[9][36] , 
        \negative_inputs[9][35] , \negative_inputs[9][34] , 
        \negative_inputs[9][33] , \negative_inputs[9][32] , 
        \negative_inputs[9][31] , \negative_inputs[9][30] , 
        \negative_inputs[9][29] , \negative_inputs[9][28] , 
        \negative_inputs[9][27] , \negative_inputs[9][26] , 
        \negative_inputs[9][25] , \negative_inputs[9][24] , 
        \negative_inputs[9][23] , \negative_inputs[9][22] , 
        \negative_inputs[9][21] , \negative_inputs[9][20] , 
        \negative_inputs[9][19] , \negative_inputs[9][18] , 
        \negative_inputs[9][17] , \negative_inputs[9][16] , 
        \negative_inputs[9][15] , \negative_inputs[9][14] , 
        \negative_inputs[9][13] , \negative_inputs[9][12] , 
        \negative_inputs[9][11] , \negative_inputs[9][10] , 
        \negative_inputs[9][9] , \negative_inputs[9][8] , 
        \negative_inputs[9][7] , \negative_inputs[9][6] , 
        \negative_inputs[9][5] , \negative_inputs[9][4] , 
        \negative_inputs[9][3] , \negative_inputs[9][2] , 
        \negative_inputs[9][1] , \negative_inputs[9][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[14:12]), .Y({\ADDER_IN_from_mux[4][63] , 
        \ADDER_IN_from_mux[4][62] , \ADDER_IN_from_mux[4][61] , 
        \ADDER_IN_from_mux[4][60] , \ADDER_IN_from_mux[4][59] , 
        \ADDER_IN_from_mux[4][58] , \ADDER_IN_from_mux[4][57] , 
        \ADDER_IN_from_mux[4][56] , \ADDER_IN_from_mux[4][55] , 
        \ADDER_IN_from_mux[4][54] , \ADDER_IN_from_mux[4][53] , 
        \ADDER_IN_from_mux[4][52] , \ADDER_IN_from_mux[4][51] , 
        \ADDER_IN_from_mux[4][50] , \ADDER_IN_from_mux[4][49] , 
        \ADDER_IN_from_mux[4][48] , \ADDER_IN_from_mux[4][47] , 
        \ADDER_IN_from_mux[4][46] , \ADDER_IN_from_mux[4][45] , 
        \ADDER_IN_from_mux[4][44] , \ADDER_IN_from_mux[4][43] , 
        \ADDER_IN_from_mux[4][42] , \ADDER_IN_from_mux[4][41] , 
        \ADDER_IN_from_mux[4][40] , \ADDER_IN_from_mux[4][39] , 
        \ADDER_IN_from_mux[4][38] , \ADDER_IN_from_mux[4][37] , 
        \ADDER_IN_from_mux[4][36] , \ADDER_IN_from_mux[4][35] , 
        \ADDER_IN_from_mux[4][34] , \ADDER_IN_from_mux[4][33] , 
        \ADDER_IN_from_mux[4][32] , \ADDER_IN_from_mux[4][31] , 
        \ADDER_IN_from_mux[4][30] , \ADDER_IN_from_mux[4][29] , 
        \ADDER_IN_from_mux[4][28] , \ADDER_IN_from_mux[4][27] , 
        \ADDER_IN_from_mux[4][26] , \ADDER_IN_from_mux[4][25] , 
        \ADDER_IN_from_mux[4][24] , \ADDER_IN_from_mux[4][23] , 
        \ADDER_IN_from_mux[4][22] , \ADDER_IN_from_mux[4][21] , 
        \ADDER_IN_from_mux[4][20] , \ADDER_IN_from_mux[4][19] , 
        \ADDER_IN_from_mux[4][18] , \ADDER_IN_from_mux[4][17] , 
        \ADDER_IN_from_mux[4][16] , \ADDER_IN_from_mux[4][15] , 
        \ADDER_IN_from_mux[4][14] , \ADDER_IN_from_mux[4][13] , 
        \ADDER_IN_from_mux[4][12] , \ADDER_IN_from_mux[4][11] , 
        \ADDER_IN_from_mux[4][10] , \ADDER_IN_from_mux[4][9] , 
        \ADDER_IN_from_mux[4][8] , \ADDER_IN_from_mux[4][7] , 
        \ADDER_IN_from_mux[4][6] , \ADDER_IN_from_mux[4][5] , 
        \ADDER_IN_from_mux[4][4] , \ADDER_IN_from_mux[4][3] , 
        \ADDER_IN_from_mux[4][2] , \ADDER_IN_from_mux[4][1] , 
        \ADDER_IN_from_mux[4][0] }) );
  MUX81_GENERIC_NBIT64_11 MUX81_N_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n665, 
        n666, n666, n666, n666, n666, n666, n666, n666, n666, n666, n666, n666, 
        n666, n666, n666, n666, n666, n666, n666, n666, n666, n666, n627, n624, 
        n618, n615, n612, n610, n606, n600, n597, n594, n588, n582, n575, n572, 
        n566, n563, n556, n553, n550, n547, n541, n538, n535, n532, n491, n527, 
        n496, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n668, n668, n668, n668, n668, n668, n668, n668, 
        n668, n668, n668, n668, n668, n668, n668, n668, n668, n668, n668, n669, 
        n669, n669, n628, n624, n619, n616, n613, n610, n606, n601, n598, n594, 
        n588, n583, n576, n572, n567, n564, n557, n554, n551, n547, n542, n537, 
        n534, n531, n491, n527, n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[10][63] , \negative_inputs[10][62] , 
        \negative_inputs[10][61] , \negative_inputs[10][60] , 
        \negative_inputs[10][59] , \negative_inputs[10][58] , 
        \negative_inputs[10][57] , \negative_inputs[10][56] , 
        \negative_inputs[10][55] , \negative_inputs[10][54] , 
        \negative_inputs[10][53] , \negative_inputs[10][52] , 
        \negative_inputs[10][51] , \negative_inputs[10][50] , 
        \negative_inputs[10][49] , \negative_inputs[10][48] , 
        \negative_inputs[10][47] , \negative_inputs[10][46] , 
        \negative_inputs[10][45] , \negative_inputs[10][44] , 
        \negative_inputs[10][43] , \negative_inputs[10][42] , 
        \negative_inputs[10][41] , \negative_inputs[10][40] , 
        \negative_inputs[10][39] , \negative_inputs[10][38] , 
        \negative_inputs[10][37] , \negative_inputs[10][36] , 
        \negative_inputs[10][35] , \negative_inputs[10][34] , 
        \negative_inputs[10][33] , \negative_inputs[10][32] , 
        \negative_inputs[10][31] , \negative_inputs[10][30] , 
        \negative_inputs[10][29] , \negative_inputs[10][28] , 
        \negative_inputs[10][27] , \negative_inputs[10][26] , 
        \negative_inputs[10][25] , \negative_inputs[10][24] , 
        \negative_inputs[10][23] , \negative_inputs[10][22] , 
        \negative_inputs[10][21] , \negative_inputs[10][20] , 
        \negative_inputs[10][19] , \negative_inputs[10][18] , 
        \negative_inputs[10][17] , \negative_inputs[10][16] , 
        \negative_inputs[10][15] , \negative_inputs[10][14] , 
        \negative_inputs[10][13] , \negative_inputs[10][12] , 
        \negative_inputs[10][11] , \negative_inputs[10][10] , 
        \negative_inputs[10][9] , \negative_inputs[10][8] , 
        \negative_inputs[10][7] , \negative_inputs[10][6] , 
        \negative_inputs[10][5] , \negative_inputs[10][4] , 
        \negative_inputs[10][3] , \negative_inputs[10][2] , 
        \negative_inputs[10][1] , \negative_inputs[10][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[11][63] , \negative_inputs[11][62] , 
        \negative_inputs[11][61] , \negative_inputs[11][60] , 
        \negative_inputs[11][59] , \negative_inputs[11][58] , 
        \negative_inputs[11][57] , \negative_inputs[11][56] , 
        \negative_inputs[11][55] , \negative_inputs[11][54] , 
        \negative_inputs[11][53] , \negative_inputs[11][52] , 
        \negative_inputs[11][51] , \negative_inputs[11][50] , 
        \negative_inputs[11][49] , \negative_inputs[11][48] , 
        \negative_inputs[11][47] , \negative_inputs[11][46] , 
        \negative_inputs[11][45] , \negative_inputs[11][44] , 
        \negative_inputs[11][43] , \negative_inputs[11][42] , 
        \negative_inputs[11][41] , \negative_inputs[11][40] , 
        \negative_inputs[11][39] , \negative_inputs[11][38] , 
        \negative_inputs[11][37] , \negative_inputs[11][36] , 
        \negative_inputs[11][35] , \negative_inputs[11][34] , 
        \negative_inputs[11][33] , \negative_inputs[11][32] , 
        \negative_inputs[11][31] , \negative_inputs[11][30] , 
        \negative_inputs[11][29] , \negative_inputs[11][28] , 
        \negative_inputs[11][27] , \negative_inputs[11][26] , 
        \negative_inputs[11][25] , \negative_inputs[11][24] , 
        \negative_inputs[11][23] , \negative_inputs[11][22] , 
        \negative_inputs[11][21] , \negative_inputs[11][20] , 
        \negative_inputs[11][19] , \negative_inputs[11][18] , 
        \negative_inputs[11][17] , \negative_inputs[11][16] , 
        \negative_inputs[11][15] , \negative_inputs[11][14] , 
        \negative_inputs[11][13] , \negative_inputs[11][12] , 
        \negative_inputs[11][11] , \negative_inputs[11][10] , 
        \negative_inputs[11][9] , \negative_inputs[11][8] , 
        \negative_inputs[11][7] , \negative_inputs[11][6] , 
        \negative_inputs[11][5] , \negative_inputs[11][4] , 
        \negative_inputs[11][3] , \negative_inputs[11][2] , 
        \negative_inputs[11][1] , \negative_inputs[11][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[17:15]), .Y({\ADDER_IN_from_mux[5][63] , 
        \ADDER_IN_from_mux[5][62] , \ADDER_IN_from_mux[5][61] , 
        \ADDER_IN_from_mux[5][60] , \ADDER_IN_from_mux[5][59] , 
        \ADDER_IN_from_mux[5][58] , \ADDER_IN_from_mux[5][57] , 
        \ADDER_IN_from_mux[5][56] , \ADDER_IN_from_mux[5][55] , 
        \ADDER_IN_from_mux[5][54] , \ADDER_IN_from_mux[5][53] , 
        \ADDER_IN_from_mux[5][52] , \ADDER_IN_from_mux[5][51] , 
        \ADDER_IN_from_mux[5][50] , \ADDER_IN_from_mux[5][49] , 
        \ADDER_IN_from_mux[5][48] , \ADDER_IN_from_mux[5][47] , 
        \ADDER_IN_from_mux[5][46] , \ADDER_IN_from_mux[5][45] , 
        \ADDER_IN_from_mux[5][44] , \ADDER_IN_from_mux[5][43] , 
        \ADDER_IN_from_mux[5][42] , \ADDER_IN_from_mux[5][41] , 
        \ADDER_IN_from_mux[5][40] , \ADDER_IN_from_mux[5][39] , 
        \ADDER_IN_from_mux[5][38] , \ADDER_IN_from_mux[5][37] , 
        \ADDER_IN_from_mux[5][36] , \ADDER_IN_from_mux[5][35] , 
        \ADDER_IN_from_mux[5][34] , \ADDER_IN_from_mux[5][33] , 
        \ADDER_IN_from_mux[5][32] , \ADDER_IN_from_mux[5][31] , 
        \ADDER_IN_from_mux[5][30] , \ADDER_IN_from_mux[5][29] , 
        \ADDER_IN_from_mux[5][28] , \ADDER_IN_from_mux[5][27] , 
        \ADDER_IN_from_mux[5][26] , \ADDER_IN_from_mux[5][25] , 
        \ADDER_IN_from_mux[5][24] , \ADDER_IN_from_mux[5][23] , 
        \ADDER_IN_from_mux[5][22] , \ADDER_IN_from_mux[5][21] , 
        \ADDER_IN_from_mux[5][20] , \ADDER_IN_from_mux[5][19] , 
        \ADDER_IN_from_mux[5][18] , \ADDER_IN_from_mux[5][17] , 
        \ADDER_IN_from_mux[5][16] , \ADDER_IN_from_mux[5][15] , 
        \ADDER_IN_from_mux[5][14] , \ADDER_IN_from_mux[5][13] , 
        \ADDER_IN_from_mux[5][12] , \ADDER_IN_from_mux[5][11] , 
        \ADDER_IN_from_mux[5][10] , \ADDER_IN_from_mux[5][9] , 
        \ADDER_IN_from_mux[5][8] , \ADDER_IN_from_mux[5][7] , 
        \ADDER_IN_from_mux[5][6] , \ADDER_IN_from_mux[5][5] , 
        \ADDER_IN_from_mux[5][4] , \ADDER_IN_from_mux[5][3] , 
        \ADDER_IN_from_mux[5][2] , \ADDER_IN_from_mux[5][1] , 
        \ADDER_IN_from_mux[5][0] }) );
  MUX81_GENERIC_NBIT64_10 MUX81_N_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n661, 
        n659, n659, n659, n660, n660, n660, n660, n660, n660, n660, n660, n660, 
        n660, n660, n660, n660, n660, n660, n660, n660, n627, n624, n619, n616, 
        n612, n610, n606, n601, n597, n594, n588, n582, n575, n572, n566, n563, 
        n556, n553, n550, n547, n541, n537, n535, n532, n530, n527, n506, n521, 
        n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n669, n669, n669, n669, n669, n669, n669, n669, 
        n669, n669, n669, n669, n669, n669, n669, n669, n669, n669, n669, n669, 
        n628, n624, n619, n616, n613, n610, n606, n601, n598, n594, n588, n583, 
        n576, n572, n567, n564, n557, n554, n551, n547, n542, n538, n535, n532, 
        n530, n527, n506, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[12][63] , \negative_inputs[12][62] , 
        \negative_inputs[12][61] , \negative_inputs[12][60] , 
        \negative_inputs[12][59] , \negative_inputs[12][58] , 
        \negative_inputs[12][57] , \negative_inputs[12][56] , 
        \negative_inputs[12][55] , \negative_inputs[12][54] , 
        \negative_inputs[12][53] , \negative_inputs[12][52] , 
        \negative_inputs[12][51] , \negative_inputs[12][50] , 
        \negative_inputs[12][49] , \negative_inputs[12][48] , 
        \negative_inputs[12][47] , \negative_inputs[12][46] , 
        \negative_inputs[12][45] , \negative_inputs[12][44] , 
        \negative_inputs[12][43] , \negative_inputs[12][42] , 
        \negative_inputs[12][41] , \negative_inputs[12][40] , 
        \negative_inputs[12][39] , \negative_inputs[12][38] , 
        \negative_inputs[12][37] , \negative_inputs[12][36] , 
        \negative_inputs[12][35] , \negative_inputs[12][34] , 
        \negative_inputs[12][33] , \negative_inputs[12][32] , 
        \negative_inputs[12][31] , \negative_inputs[12][30] , 
        \negative_inputs[12][29] , \negative_inputs[12][28] , 
        \negative_inputs[12][27] , \negative_inputs[12][26] , 
        \negative_inputs[12][25] , \negative_inputs[12][24] , 
        \negative_inputs[12][23] , \negative_inputs[12][22] , 
        \negative_inputs[12][21] , \negative_inputs[12][20] , 
        \negative_inputs[12][19] , \negative_inputs[12][18] , 
        \negative_inputs[12][17] , \negative_inputs[12][16] , 
        \negative_inputs[12][15] , \negative_inputs[12][14] , 
        \negative_inputs[12][13] , \negative_inputs[12][12] , 
        \negative_inputs[12][11] , \negative_inputs[12][10] , 
        \negative_inputs[12][9] , \negative_inputs[12][8] , 
        \negative_inputs[12][7] , \negative_inputs[12][6] , 
        \negative_inputs[12][5] , \negative_inputs[12][4] , 
        \negative_inputs[12][3] , \negative_inputs[12][2] , 
        \negative_inputs[12][1] , \negative_inputs[12][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[13][63] , \negative_inputs[13][62] , 
        \negative_inputs[13][61] , \negative_inputs[13][60] , 
        \negative_inputs[13][59] , \negative_inputs[13][58] , 
        \negative_inputs[13][57] , \negative_inputs[13][56] , 
        \negative_inputs[13][55] , \negative_inputs[13][54] , 
        \negative_inputs[13][53] , \negative_inputs[13][52] , 
        \negative_inputs[13][51] , \negative_inputs[13][50] , 
        \negative_inputs[13][49] , \negative_inputs[13][48] , 
        \negative_inputs[13][47] , \negative_inputs[13][46] , 
        \negative_inputs[13][45] , \negative_inputs[13][44] , 
        \negative_inputs[13][43] , \negative_inputs[13][42] , 
        \negative_inputs[13][41] , \negative_inputs[13][40] , 
        \negative_inputs[13][39] , \negative_inputs[13][38] , 
        \negative_inputs[13][37] , \negative_inputs[13][36] , 
        \negative_inputs[13][35] , \negative_inputs[13][34] , 
        \negative_inputs[13][33] , \negative_inputs[13][32] , 
        \negative_inputs[13][31] , \negative_inputs[13][30] , 
        \negative_inputs[13][29] , \negative_inputs[13][28] , 
        \negative_inputs[13][27] , \negative_inputs[13][26] , 
        \negative_inputs[13][25] , \negative_inputs[13][24] , 
        \negative_inputs[13][23] , \negative_inputs[13][22] , 
        \negative_inputs[13][21] , \negative_inputs[13][20] , 
        \negative_inputs[13][19] , \negative_inputs[13][18] , 
        \negative_inputs[13][17] , \negative_inputs[13][16] , 
        \negative_inputs[13][15] , \negative_inputs[13][14] , 
        \negative_inputs[13][13] , \negative_inputs[13][12] , 
        \negative_inputs[13][11] , \negative_inputs[13][10] , 
        \negative_inputs[13][9] , \negative_inputs[13][8] , 
        \negative_inputs[13][7] , \negative_inputs[13][6] , 
        \negative_inputs[13][5] , \negative_inputs[13][4] , 
        \negative_inputs[13][3] , \negative_inputs[13][2] , 
        \negative_inputs[13][1] , \negative_inputs[13][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[20:18]), .Y({\ADDER_IN_from_mux[6][63] , 
        \ADDER_IN_from_mux[6][62] , \ADDER_IN_from_mux[6][61] , 
        \ADDER_IN_from_mux[6][60] , \ADDER_IN_from_mux[6][59] , 
        \ADDER_IN_from_mux[6][58] , \ADDER_IN_from_mux[6][57] , 
        \ADDER_IN_from_mux[6][56] , \ADDER_IN_from_mux[6][55] , 
        \ADDER_IN_from_mux[6][54] , \ADDER_IN_from_mux[6][53] , 
        \ADDER_IN_from_mux[6][52] , \ADDER_IN_from_mux[6][51] , 
        \ADDER_IN_from_mux[6][50] , \ADDER_IN_from_mux[6][49] , 
        \ADDER_IN_from_mux[6][48] , \ADDER_IN_from_mux[6][47] , 
        \ADDER_IN_from_mux[6][46] , \ADDER_IN_from_mux[6][45] , 
        \ADDER_IN_from_mux[6][44] , \ADDER_IN_from_mux[6][43] , 
        \ADDER_IN_from_mux[6][42] , \ADDER_IN_from_mux[6][41] , 
        \ADDER_IN_from_mux[6][40] , \ADDER_IN_from_mux[6][39] , 
        \ADDER_IN_from_mux[6][38] , \ADDER_IN_from_mux[6][37] , 
        \ADDER_IN_from_mux[6][36] , \ADDER_IN_from_mux[6][35] , 
        \ADDER_IN_from_mux[6][34] , \ADDER_IN_from_mux[6][33] , 
        \ADDER_IN_from_mux[6][32] , \ADDER_IN_from_mux[6][31] , 
        \ADDER_IN_from_mux[6][30] , \ADDER_IN_from_mux[6][29] , 
        \ADDER_IN_from_mux[6][28] , \ADDER_IN_from_mux[6][27] , 
        \ADDER_IN_from_mux[6][26] , \ADDER_IN_from_mux[6][25] , 
        \ADDER_IN_from_mux[6][24] , \ADDER_IN_from_mux[6][23] , 
        \ADDER_IN_from_mux[6][22] , \ADDER_IN_from_mux[6][21] , 
        \ADDER_IN_from_mux[6][20] , \ADDER_IN_from_mux[6][19] , 
        \ADDER_IN_from_mux[6][18] , \ADDER_IN_from_mux[6][17] , 
        \ADDER_IN_from_mux[6][16] , \ADDER_IN_from_mux[6][15] , 
        \ADDER_IN_from_mux[6][14] , \ADDER_IN_from_mux[6][13] , 
        \ADDER_IN_from_mux[6][12] , \ADDER_IN_from_mux[6][11] , 
        \ADDER_IN_from_mux[6][10] , \ADDER_IN_from_mux[6][9] , 
        \ADDER_IN_from_mux[6][8] , \ADDER_IN_from_mux[6][7] , 
        \ADDER_IN_from_mux[6][6] , \ADDER_IN_from_mux[6][5] , 
        \ADDER_IN_from_mux[6][4] , \ADDER_IN_from_mux[6][3] , 
        \ADDER_IN_from_mux[6][2] , \ADDER_IN_from_mux[6][1] , 
        \ADDER_IN_from_mux[6][0] }) );
  MUX81_GENERIC_NBIT64_9 MUX81_N_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n660, 
        n660, n660, n660, n660, n660, n660, n660, n660, n660, n660, n660, n660, 
        n660, n660, n660, n660, n660, n659, n627, n624, n619, n616, n612, n609, 
        n606, n601, n597, n594, n588, n582, n575, n572, n567, n563, n556, n553, 
        n550, n547, n541, n537, n535, n531, n530, n527, n496, n521, n517, n515, 
        n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n670, n670, n670, n670, n670, n670, n670, n670, 
        n670, n670, n670, n670, n670, n670, n670, n670, n670, n670, n628, n624, 
        n619, n616, n613, n610, n606, n601, n598, n594, n588, n583, n576, n572, 
        n567, n564, n557, n554, n551, n547, n542, n537, n535, n531, n530, n527, 
        n506, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[14][63] , \negative_inputs[14][62] , 
        \negative_inputs[14][61] , \negative_inputs[14][60] , 
        \negative_inputs[14][59] , \negative_inputs[14][58] , 
        \negative_inputs[14][57] , \negative_inputs[14][56] , 
        \negative_inputs[14][55] , \negative_inputs[14][54] , 
        \negative_inputs[14][53] , \negative_inputs[14][52] , 
        \negative_inputs[14][51] , \negative_inputs[14][50] , 
        \negative_inputs[14][49] , \negative_inputs[14][48] , 
        \negative_inputs[14][47] , \negative_inputs[14][46] , 
        \negative_inputs[14][45] , \negative_inputs[14][44] , 
        \negative_inputs[14][43] , \negative_inputs[14][42] , 
        \negative_inputs[14][41] , \negative_inputs[14][40] , 
        \negative_inputs[14][39] , \negative_inputs[14][38] , 
        \negative_inputs[14][37] , \negative_inputs[14][36] , 
        \negative_inputs[14][35] , \negative_inputs[14][34] , 
        \negative_inputs[14][33] , \negative_inputs[14][32] , 
        \negative_inputs[14][31] , \negative_inputs[14][30] , 
        \negative_inputs[14][29] , \negative_inputs[14][28] , 
        \negative_inputs[14][27] , \negative_inputs[14][26] , 
        \negative_inputs[14][25] , \negative_inputs[14][24] , 
        \negative_inputs[14][23] , \negative_inputs[14][22] , 
        \negative_inputs[14][21] , \negative_inputs[14][20] , 
        \negative_inputs[14][19] , \negative_inputs[14][18] , 
        \negative_inputs[14][17] , \negative_inputs[14][16] , 
        \negative_inputs[14][15] , \negative_inputs[14][14] , 
        \negative_inputs[14][13] , \negative_inputs[14][12] , 
        \negative_inputs[14][11] , \negative_inputs[14][10] , 
        \negative_inputs[14][9] , \negative_inputs[14][8] , 
        \negative_inputs[14][7] , \negative_inputs[14][6] , 
        \negative_inputs[14][5] , \negative_inputs[14][4] , 
        \negative_inputs[14][3] , \negative_inputs[14][2] , 
        \negative_inputs[14][1] , \negative_inputs[14][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[15][63] , \negative_inputs[15][62] , 
        \negative_inputs[15][61] , \negative_inputs[15][60] , 
        \negative_inputs[15][59] , \negative_inputs[15][58] , 
        \negative_inputs[15][57] , \negative_inputs[15][56] , 
        \negative_inputs[15][55] , \negative_inputs[15][54] , 
        \negative_inputs[15][53] , \negative_inputs[15][52] , 
        \negative_inputs[15][51] , \negative_inputs[15][50] , 
        \negative_inputs[15][49] , \negative_inputs[15][48] , 
        \negative_inputs[15][47] , \negative_inputs[15][46] , 
        \negative_inputs[15][45] , \negative_inputs[15][44] , 
        \negative_inputs[15][43] , \negative_inputs[15][42] , 
        \negative_inputs[15][41] , \negative_inputs[15][40] , 
        \negative_inputs[15][39] , \negative_inputs[15][38] , 
        \negative_inputs[15][37] , \negative_inputs[15][36] , 
        \negative_inputs[15][35] , \negative_inputs[15][34] , 
        \negative_inputs[15][33] , \negative_inputs[15][32] , 
        \negative_inputs[15][31] , \negative_inputs[15][30] , 
        \negative_inputs[15][29] , \negative_inputs[15][28] , 
        \negative_inputs[15][27] , \negative_inputs[15][26] , 
        \negative_inputs[15][25] , \negative_inputs[15][24] , 
        \negative_inputs[15][23] , \negative_inputs[15][22] , 
        \negative_inputs[15][21] , \negative_inputs[15][20] , 
        \negative_inputs[15][19] , \negative_inputs[15][18] , 
        \negative_inputs[15][17] , \negative_inputs[15][16] , 
        \negative_inputs[15][15] , \negative_inputs[15][14] , 
        \negative_inputs[15][13] , \negative_inputs[15][12] , 
        \negative_inputs[15][11] , \negative_inputs[15][10] , 
        \negative_inputs[15][9] , \negative_inputs[15][8] , 
        \negative_inputs[15][7] , \negative_inputs[15][6] , 
        \negative_inputs[15][5] , \negative_inputs[15][4] , 
        \negative_inputs[15][3] , \negative_inputs[15][2] , 
        \negative_inputs[15][1] , \negative_inputs[15][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[23:21]), .Y({\ADDER_IN_from_mux[7][63] , 
        \ADDER_IN_from_mux[7][62] , \ADDER_IN_from_mux[7][61] , 
        \ADDER_IN_from_mux[7][60] , \ADDER_IN_from_mux[7][59] , 
        \ADDER_IN_from_mux[7][58] , \ADDER_IN_from_mux[7][57] , 
        \ADDER_IN_from_mux[7][56] , \ADDER_IN_from_mux[7][55] , 
        \ADDER_IN_from_mux[7][54] , \ADDER_IN_from_mux[7][53] , 
        \ADDER_IN_from_mux[7][52] , \ADDER_IN_from_mux[7][51] , 
        \ADDER_IN_from_mux[7][50] , \ADDER_IN_from_mux[7][49] , 
        \ADDER_IN_from_mux[7][48] , \ADDER_IN_from_mux[7][47] , 
        \ADDER_IN_from_mux[7][46] , \ADDER_IN_from_mux[7][45] , 
        \ADDER_IN_from_mux[7][44] , \ADDER_IN_from_mux[7][43] , 
        \ADDER_IN_from_mux[7][42] , \ADDER_IN_from_mux[7][41] , 
        \ADDER_IN_from_mux[7][40] , \ADDER_IN_from_mux[7][39] , 
        \ADDER_IN_from_mux[7][38] , \ADDER_IN_from_mux[7][37] , 
        \ADDER_IN_from_mux[7][36] , \ADDER_IN_from_mux[7][35] , 
        \ADDER_IN_from_mux[7][34] , \ADDER_IN_from_mux[7][33] , 
        \ADDER_IN_from_mux[7][32] , \ADDER_IN_from_mux[7][31] , 
        \ADDER_IN_from_mux[7][30] , \ADDER_IN_from_mux[7][29] , 
        \ADDER_IN_from_mux[7][28] , \ADDER_IN_from_mux[7][27] , 
        \ADDER_IN_from_mux[7][26] , \ADDER_IN_from_mux[7][25] , 
        \ADDER_IN_from_mux[7][24] , \ADDER_IN_from_mux[7][23] , 
        \ADDER_IN_from_mux[7][22] , \ADDER_IN_from_mux[7][21] , 
        \ADDER_IN_from_mux[7][20] , \ADDER_IN_from_mux[7][19] , 
        \ADDER_IN_from_mux[7][18] , \ADDER_IN_from_mux[7][17] , 
        \ADDER_IN_from_mux[7][16] , \ADDER_IN_from_mux[7][15] , 
        \ADDER_IN_from_mux[7][14] , \ADDER_IN_from_mux[7][13] , 
        \ADDER_IN_from_mux[7][12] , \ADDER_IN_from_mux[7][11] , 
        \ADDER_IN_from_mux[7][10] , \ADDER_IN_from_mux[7][9] , 
        \ADDER_IN_from_mux[7][8] , \ADDER_IN_from_mux[7][7] , 
        \ADDER_IN_from_mux[7][6] , \ADDER_IN_from_mux[7][5] , 
        \ADDER_IN_from_mux[7][4] , \ADDER_IN_from_mux[7][3] , 
        \ADDER_IN_from_mux[7][2] , \ADDER_IN_from_mux[7][1] , 
        \ADDER_IN_from_mux[7][0] }) );
  MUX81_GENERIC_NBIT64_8 MUX81_N_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n661, 
        n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, 
        n661, n661, n661, n661, n627, n624, n619, n616, n612, n610, n606, n601, 
        n598, n594, n588, n582, n575, n572, n566, n563, n556, n553, n551, n547, 
        n541, n538, n535, n532, n491, n527, n506, n521, n517, n515, n507, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n670, n670, n670, n670, n669, n669, n669, n669, 
        n669, n669, n669, n669, n669, n669, n669, n669, n628, n625, n619, n616, 
        n613, n610, n606, n601, n598, n594, n588, n583, n576, n572, n567, n564, 
        n557, n554, n551, n547, n542, n537, n534, n532, n530, n527, n506, n521, 
        n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[16][63] , \negative_inputs[16][62] , 
        \negative_inputs[16][61] , \negative_inputs[16][60] , 
        \negative_inputs[16][59] , \negative_inputs[16][58] , 
        \negative_inputs[16][57] , \negative_inputs[16][56] , 
        \negative_inputs[16][55] , \negative_inputs[16][54] , 
        \negative_inputs[16][53] , \negative_inputs[16][52] , 
        \negative_inputs[16][51] , \negative_inputs[16][50] , 
        \negative_inputs[16][49] , \negative_inputs[16][48] , 
        \negative_inputs[16][47] , \negative_inputs[16][46] , 
        \negative_inputs[16][45] , \negative_inputs[16][44] , 
        \negative_inputs[16][43] , \negative_inputs[16][42] , 
        \negative_inputs[16][41] , \negative_inputs[16][40] , 
        \negative_inputs[16][39] , \negative_inputs[16][38] , 
        \negative_inputs[16][37] , \negative_inputs[16][36] , 
        \negative_inputs[16][35] , \negative_inputs[16][34] , 
        \negative_inputs[16][33] , \negative_inputs[16][32] , 
        \negative_inputs[16][31] , \negative_inputs[16][30] , 
        \negative_inputs[16][29] , \negative_inputs[16][28] , 
        \negative_inputs[16][27] , \negative_inputs[16][26] , 
        \negative_inputs[16][25] , \negative_inputs[16][24] , 
        \negative_inputs[16][23] , \negative_inputs[16][22] , 
        \negative_inputs[16][21] , \negative_inputs[16][20] , 
        \negative_inputs[16][19] , \negative_inputs[16][18] , 
        \negative_inputs[16][17] , \negative_inputs[16][16] , 
        \negative_inputs[16][15] , \negative_inputs[16][14] , 
        \negative_inputs[16][13] , \negative_inputs[16][12] , 
        \negative_inputs[16][11] , \negative_inputs[16][10] , 
        \negative_inputs[16][9] , \negative_inputs[16][8] , 
        \negative_inputs[16][7] , \negative_inputs[16][6] , 
        \negative_inputs[16][5] , \negative_inputs[16][4] , 
        \negative_inputs[16][3] , \negative_inputs[16][2] , 
        \negative_inputs[16][1] , \negative_inputs[16][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[17][63] , \negative_inputs[17][62] , 
        \negative_inputs[17][61] , \negative_inputs[17][60] , 
        \negative_inputs[17][59] , \negative_inputs[17][58] , 
        \negative_inputs[17][57] , \negative_inputs[17][56] , 
        \negative_inputs[17][55] , \negative_inputs[17][54] , 
        \negative_inputs[17][53] , \negative_inputs[17][52] , 
        \negative_inputs[17][51] , \negative_inputs[17][50] , 
        \negative_inputs[17][49] , \negative_inputs[17][48] , 
        \negative_inputs[17][47] , \negative_inputs[17][46] , 
        \negative_inputs[17][45] , \negative_inputs[17][44] , 
        \negative_inputs[17][43] , \negative_inputs[17][42] , 
        \negative_inputs[17][41] , \negative_inputs[17][40] , 
        \negative_inputs[17][39] , \negative_inputs[17][38] , 
        \negative_inputs[17][37] , \negative_inputs[17][36] , 
        \negative_inputs[17][35] , \negative_inputs[17][34] , 
        \negative_inputs[17][33] , \negative_inputs[17][32] , 
        \negative_inputs[17][31] , \negative_inputs[17][30] , 
        \negative_inputs[17][29] , \negative_inputs[17][28] , 
        \negative_inputs[17][27] , \negative_inputs[17][26] , 
        \negative_inputs[17][25] , \negative_inputs[17][24] , 
        \negative_inputs[17][23] , \negative_inputs[17][22] , 
        \negative_inputs[17][21] , \negative_inputs[17][20] , 
        \negative_inputs[17][19] , \negative_inputs[17][18] , 
        \negative_inputs[17][17] , \negative_inputs[17][16] , 
        \negative_inputs[17][15] , \negative_inputs[17][14] , 
        \negative_inputs[17][13] , \negative_inputs[17][12] , 
        \negative_inputs[17][11] , \negative_inputs[17][10] , 
        \negative_inputs[17][9] , \negative_inputs[17][8] , 
        \negative_inputs[17][7] , \negative_inputs[17][6] , 
        \negative_inputs[17][5] , \negative_inputs[17][4] , 
        \negative_inputs[17][3] , \negative_inputs[17][2] , 
        \negative_inputs[17][1] , \negative_inputs[17][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[26:24]), .Y({\ADDER_IN_from_mux[8][63] , 
        \ADDER_IN_from_mux[8][62] , \ADDER_IN_from_mux[8][61] , 
        \ADDER_IN_from_mux[8][60] , \ADDER_IN_from_mux[8][59] , 
        \ADDER_IN_from_mux[8][58] , \ADDER_IN_from_mux[8][57] , 
        \ADDER_IN_from_mux[8][56] , \ADDER_IN_from_mux[8][55] , 
        \ADDER_IN_from_mux[8][54] , \ADDER_IN_from_mux[8][53] , 
        \ADDER_IN_from_mux[8][52] , \ADDER_IN_from_mux[8][51] , 
        \ADDER_IN_from_mux[8][50] , \ADDER_IN_from_mux[8][49] , 
        \ADDER_IN_from_mux[8][48] , \ADDER_IN_from_mux[8][47] , 
        \ADDER_IN_from_mux[8][46] , \ADDER_IN_from_mux[8][45] , 
        \ADDER_IN_from_mux[8][44] , \ADDER_IN_from_mux[8][43] , 
        \ADDER_IN_from_mux[8][42] , \ADDER_IN_from_mux[8][41] , 
        \ADDER_IN_from_mux[8][40] , \ADDER_IN_from_mux[8][39] , 
        \ADDER_IN_from_mux[8][38] , \ADDER_IN_from_mux[8][37] , 
        \ADDER_IN_from_mux[8][36] , \ADDER_IN_from_mux[8][35] , 
        \ADDER_IN_from_mux[8][34] , \ADDER_IN_from_mux[8][33] , 
        \ADDER_IN_from_mux[8][32] , \ADDER_IN_from_mux[8][31] , 
        \ADDER_IN_from_mux[8][30] , \ADDER_IN_from_mux[8][29] , 
        \ADDER_IN_from_mux[8][28] , \ADDER_IN_from_mux[8][27] , 
        \ADDER_IN_from_mux[8][26] , \ADDER_IN_from_mux[8][25] , 
        \ADDER_IN_from_mux[8][24] , \ADDER_IN_from_mux[8][23] , 
        \ADDER_IN_from_mux[8][22] , \ADDER_IN_from_mux[8][21] , 
        \ADDER_IN_from_mux[8][20] , \ADDER_IN_from_mux[8][19] , 
        \ADDER_IN_from_mux[8][18] , \ADDER_IN_from_mux[8][17] , 
        \ADDER_IN_from_mux[8][16] , \ADDER_IN_from_mux[8][15] , 
        \ADDER_IN_from_mux[8][14] , \ADDER_IN_from_mux[8][13] , 
        \ADDER_IN_from_mux[8][12] , \ADDER_IN_from_mux[8][11] , 
        \ADDER_IN_from_mux[8][10] , \ADDER_IN_from_mux[8][9] , 
        \ADDER_IN_from_mux[8][8] , \ADDER_IN_from_mux[8][7] , 
        \ADDER_IN_from_mux[8][6] , \ADDER_IN_from_mux[8][5] , 
        \ADDER_IN_from_mux[8][4] , \ADDER_IN_from_mux[8][3] , 
        \ADDER_IN_from_mux[8][2] , \ADDER_IN_from_mux[8][1] , 
        \ADDER_IN_from_mux[8][0] }) );
  MUX81_GENERIC_NBIT64_7 MUX81_N_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n661, 
        n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, n661, 
        n661, n661, n627, n624, n619, n616, n612, n610, n606, n601, n598, n594, 
        n588, n582, n576, n572, n567, n563, n557, n553, n551, n547, n542, n537, 
        n535, n531, n530, n527, n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n669, n668, n668, n668, n668, n668, n667, n667, 
        n667, n667, n667, n667, n667, n667, n628, n625, n619, n616, n613, n610, 
        n606, n601, n598, n594, n588, n583, n576, n572, n567, n564, n557, n554, 
        n551, n547, n542, n538, n534, n531, n491, n527, n506, n521, n517, n515, 
        n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[18][63] , \negative_inputs[18][62] , 
        \negative_inputs[18][61] , \negative_inputs[18][60] , 
        \negative_inputs[18][59] , \negative_inputs[18][58] , 
        \negative_inputs[18][57] , \negative_inputs[18][56] , 
        \negative_inputs[18][55] , \negative_inputs[18][54] , 
        \negative_inputs[18][53] , \negative_inputs[18][52] , 
        \negative_inputs[18][51] , \negative_inputs[18][50] , 
        \negative_inputs[18][49] , \negative_inputs[18][48] , 
        \negative_inputs[18][47] , \negative_inputs[18][46] , 
        \negative_inputs[18][45] , \negative_inputs[18][44] , 
        \negative_inputs[18][43] , \negative_inputs[18][42] , 
        \negative_inputs[18][41] , \negative_inputs[18][40] , 
        \negative_inputs[18][39] , \negative_inputs[18][38] , 
        \negative_inputs[18][37] , \negative_inputs[18][36] , 
        \negative_inputs[18][35] , \negative_inputs[18][34] , 
        \negative_inputs[18][33] , \negative_inputs[18][32] , 
        \negative_inputs[18][31] , \negative_inputs[18][30] , 
        \negative_inputs[18][29] , \negative_inputs[18][28] , 
        \negative_inputs[18][27] , \negative_inputs[18][26] , 
        \negative_inputs[18][25] , \negative_inputs[18][24] , 
        \negative_inputs[18][23] , \negative_inputs[18][22] , 
        \negative_inputs[18][21] , \negative_inputs[18][20] , 
        \negative_inputs[18][19] , \negative_inputs[18][18] , 
        \negative_inputs[18][17] , \negative_inputs[18][16] , 
        \negative_inputs[18][15] , \negative_inputs[18][14] , 
        \negative_inputs[18][13] , \negative_inputs[18][12] , 
        \negative_inputs[18][11] , \negative_inputs[18][10] , 
        \negative_inputs[18][9] , \negative_inputs[18][8] , 
        \negative_inputs[18][7] , \negative_inputs[18][6] , 
        \negative_inputs[18][5] , \negative_inputs[18][4] , 
        \negative_inputs[18][3] , \negative_inputs[18][2] , 
        \negative_inputs[18][1] , \negative_inputs[18][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[19][63] , \negative_inputs[19][62] , 
        \negative_inputs[19][61] , \negative_inputs[19][60] , 
        \negative_inputs[19][59] , \negative_inputs[19][58] , 
        \negative_inputs[19][57] , \negative_inputs[19][56] , 
        \negative_inputs[19][55] , \negative_inputs[19][54] , 
        \negative_inputs[19][53] , \negative_inputs[19][52] , 
        \negative_inputs[19][51] , \negative_inputs[19][50] , 
        \negative_inputs[19][49] , \negative_inputs[19][48] , 
        \negative_inputs[19][47] , \negative_inputs[19][46] , 
        \negative_inputs[19][45] , \negative_inputs[19][44] , 
        \negative_inputs[19][43] , \negative_inputs[19][42] , 
        \negative_inputs[19][41] , \negative_inputs[19][40] , 
        \negative_inputs[19][39] , \negative_inputs[19][38] , 
        \negative_inputs[19][37] , \negative_inputs[19][36] , 
        \negative_inputs[19][35] , \negative_inputs[19][34] , 
        \negative_inputs[19][33] , \negative_inputs[19][32] , 
        \negative_inputs[19][31] , \negative_inputs[19][30] , 
        \negative_inputs[19][29] , \negative_inputs[19][28] , 
        \negative_inputs[19][27] , \negative_inputs[19][26] , 
        \negative_inputs[19][25] , \negative_inputs[19][24] , 
        \negative_inputs[19][23] , \negative_inputs[19][22] , 
        \negative_inputs[19][21] , \negative_inputs[19][20] , 
        \negative_inputs[19][19] , \negative_inputs[19][18] , 
        \negative_inputs[19][17] , \negative_inputs[19][16] , 
        \negative_inputs[19][15] , \negative_inputs[19][14] , 
        \negative_inputs[19][13] , \negative_inputs[19][12] , 
        \negative_inputs[19][11] , \negative_inputs[19][10] , 
        \negative_inputs[19][9] , \negative_inputs[19][8] , 
        \negative_inputs[19][7] , \negative_inputs[19][6] , 
        \negative_inputs[19][5] , \negative_inputs[19][4] , 
        \negative_inputs[19][3] , \negative_inputs[19][2] , 
        \negative_inputs[19][1] , \negative_inputs[19][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[29:27]), .Y({\ADDER_IN_from_mux[9][63] , 
        \ADDER_IN_from_mux[9][62] , \ADDER_IN_from_mux[9][61] , 
        \ADDER_IN_from_mux[9][60] , \ADDER_IN_from_mux[9][59] , 
        \ADDER_IN_from_mux[9][58] , \ADDER_IN_from_mux[9][57] , 
        \ADDER_IN_from_mux[9][56] , \ADDER_IN_from_mux[9][55] , 
        \ADDER_IN_from_mux[9][54] , \ADDER_IN_from_mux[9][53] , 
        \ADDER_IN_from_mux[9][52] , \ADDER_IN_from_mux[9][51] , 
        \ADDER_IN_from_mux[9][50] , \ADDER_IN_from_mux[9][49] , 
        \ADDER_IN_from_mux[9][48] , \ADDER_IN_from_mux[9][47] , 
        \ADDER_IN_from_mux[9][46] , \ADDER_IN_from_mux[9][45] , 
        \ADDER_IN_from_mux[9][44] , \ADDER_IN_from_mux[9][43] , 
        \ADDER_IN_from_mux[9][42] , \ADDER_IN_from_mux[9][41] , 
        \ADDER_IN_from_mux[9][40] , \ADDER_IN_from_mux[9][39] , 
        \ADDER_IN_from_mux[9][38] , \ADDER_IN_from_mux[9][37] , 
        \ADDER_IN_from_mux[9][36] , \ADDER_IN_from_mux[9][35] , 
        \ADDER_IN_from_mux[9][34] , \ADDER_IN_from_mux[9][33] , 
        \ADDER_IN_from_mux[9][32] , \ADDER_IN_from_mux[9][31] , 
        \ADDER_IN_from_mux[9][30] , \ADDER_IN_from_mux[9][29] , 
        \ADDER_IN_from_mux[9][28] , \ADDER_IN_from_mux[9][27] , 
        \ADDER_IN_from_mux[9][26] , \ADDER_IN_from_mux[9][25] , 
        \ADDER_IN_from_mux[9][24] , \ADDER_IN_from_mux[9][23] , 
        \ADDER_IN_from_mux[9][22] , \ADDER_IN_from_mux[9][21] , 
        \ADDER_IN_from_mux[9][20] , \ADDER_IN_from_mux[9][19] , 
        \ADDER_IN_from_mux[9][18] , \ADDER_IN_from_mux[9][17] , 
        \ADDER_IN_from_mux[9][16] , \ADDER_IN_from_mux[9][15] , 
        \ADDER_IN_from_mux[9][14] , \ADDER_IN_from_mux[9][13] , 
        \ADDER_IN_from_mux[9][12] , \ADDER_IN_from_mux[9][11] , 
        \ADDER_IN_from_mux[9][10] , \ADDER_IN_from_mux[9][9] , 
        \ADDER_IN_from_mux[9][8] , \ADDER_IN_from_mux[9][7] , 
        \ADDER_IN_from_mux[9][6] , \ADDER_IN_from_mux[9][5] , 
        \ADDER_IN_from_mux[9][4] , \ADDER_IN_from_mux[9][3] , 
        \ADDER_IN_from_mux[9][2] , \ADDER_IN_from_mux[9][1] , 
        \ADDER_IN_from_mux[9][0] }) );
  MUX81_GENERIC_NBIT64_6 MUX81_N_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n661, 
        n661, n662, n662, n662, n662, n662, n662, n662, n662, n662, n662, n662, 
        n627, n624, n619, n616, n612, n610, n606, n601, n598, n594, n588, n582, 
        n576, n572, n567, n563, n557, n553, n551, n547, n542, n538, n535, n532, 
        n530, n527, n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n667, n667, n666, n666, n666, n666, n666, n666, 
        n666, n668, n673, n672, n628, n625, n619, n616, n613, n610, n606, n601, 
        n598, n594, n588, n583, n576, n572, n567, n564, n557, n554, n551, n547, 
        n542, n537, n535, n531, n530, n527, n506, n521, n517, n515, n507, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[20][63] , \negative_inputs[20][62] , 
        \negative_inputs[20][61] , \negative_inputs[20][60] , 
        \negative_inputs[20][59] , \negative_inputs[20][58] , 
        \negative_inputs[20][57] , \negative_inputs[20][56] , 
        \negative_inputs[20][55] , \negative_inputs[20][54] , 
        \negative_inputs[20][53] , \negative_inputs[20][52] , 
        \negative_inputs[20][51] , \negative_inputs[20][50] , 
        \negative_inputs[20][49] , \negative_inputs[20][48] , 
        \negative_inputs[20][47] , \negative_inputs[20][46] , 
        \negative_inputs[20][45] , \negative_inputs[20][44] , 
        \negative_inputs[20][43] , \negative_inputs[20][42] , 
        \negative_inputs[20][41] , \negative_inputs[20][40] , 
        \negative_inputs[20][39] , \negative_inputs[20][38] , 
        \negative_inputs[20][37] , \negative_inputs[20][36] , 
        \negative_inputs[20][35] , \negative_inputs[20][34] , 
        \negative_inputs[20][33] , \negative_inputs[20][32] , 
        \negative_inputs[20][31] , \negative_inputs[20][30] , 
        \negative_inputs[20][29] , \negative_inputs[20][28] , 
        \negative_inputs[20][27] , \negative_inputs[20][26] , 
        \negative_inputs[20][25] , \negative_inputs[20][24] , 
        \negative_inputs[20][23] , \negative_inputs[20][22] , 
        \negative_inputs[20][21] , \negative_inputs[20][20] , 
        \negative_inputs[20][19] , \negative_inputs[20][18] , 
        \negative_inputs[20][17] , \negative_inputs[20][16] , 
        \negative_inputs[20][15] , \negative_inputs[20][14] , 
        \negative_inputs[20][13] , \negative_inputs[20][12] , 
        \negative_inputs[20][11] , \negative_inputs[20][10] , 
        \negative_inputs[20][9] , \negative_inputs[20][8] , 
        \negative_inputs[20][7] , \negative_inputs[20][6] , 
        \negative_inputs[20][5] , \negative_inputs[20][4] , 
        \negative_inputs[20][3] , \negative_inputs[20][2] , 
        \negative_inputs[20][1] , \negative_inputs[20][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[21][63] , \negative_inputs[21][62] , 
        \negative_inputs[21][61] , \negative_inputs[21][60] , 
        \negative_inputs[21][59] , \negative_inputs[21][58] , 
        \negative_inputs[21][57] , \negative_inputs[21][56] , 
        \negative_inputs[21][55] , \negative_inputs[21][54] , 
        \negative_inputs[21][53] , \negative_inputs[21][52] , 
        \negative_inputs[21][51] , \negative_inputs[21][50] , 
        \negative_inputs[21][49] , \negative_inputs[21][48] , 
        \negative_inputs[21][47] , \negative_inputs[21][46] , 
        \negative_inputs[21][45] , \negative_inputs[21][44] , 
        \negative_inputs[21][43] , \negative_inputs[21][42] , 
        \negative_inputs[21][41] , \negative_inputs[21][40] , 
        \negative_inputs[21][39] , \negative_inputs[21][38] , 
        \negative_inputs[21][37] , \negative_inputs[21][36] , 
        \negative_inputs[21][35] , \negative_inputs[21][34] , 
        \negative_inputs[21][33] , \negative_inputs[21][32] , 
        \negative_inputs[21][31] , \negative_inputs[21][30] , 
        \negative_inputs[21][29] , \negative_inputs[21][28] , 
        \negative_inputs[21][27] , \negative_inputs[21][26] , 
        \negative_inputs[21][25] , \negative_inputs[21][24] , 
        \negative_inputs[21][23] , \negative_inputs[21][22] , 
        \negative_inputs[21][21] , \negative_inputs[21][20] , 
        \negative_inputs[21][19] , \negative_inputs[21][18] , 
        \negative_inputs[21][17] , \negative_inputs[21][16] , 
        \negative_inputs[21][15] , \negative_inputs[21][14] , 
        \negative_inputs[21][13] , \negative_inputs[21][12] , 
        \negative_inputs[21][11] , \negative_inputs[21][10] , 
        \negative_inputs[21][9] , \negative_inputs[21][8] , 
        \negative_inputs[21][7] , \negative_inputs[21][6] , 
        \negative_inputs[21][5] , \negative_inputs[21][4] , 
        \negative_inputs[21][3] , \negative_inputs[21][2] , 
        \negative_inputs[21][1] , \negative_inputs[21][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[32:30]), .Y({
        \ADDER_IN_from_mux[10][63] , \ADDER_IN_from_mux[10][62] , 
        \ADDER_IN_from_mux[10][61] , \ADDER_IN_from_mux[10][60] , 
        \ADDER_IN_from_mux[10][59] , \ADDER_IN_from_mux[10][58] , 
        \ADDER_IN_from_mux[10][57] , \ADDER_IN_from_mux[10][56] , 
        \ADDER_IN_from_mux[10][55] , \ADDER_IN_from_mux[10][54] , 
        \ADDER_IN_from_mux[10][53] , \ADDER_IN_from_mux[10][52] , 
        \ADDER_IN_from_mux[10][51] , \ADDER_IN_from_mux[10][50] , 
        \ADDER_IN_from_mux[10][49] , \ADDER_IN_from_mux[10][48] , 
        \ADDER_IN_from_mux[10][47] , \ADDER_IN_from_mux[10][46] , 
        \ADDER_IN_from_mux[10][45] , \ADDER_IN_from_mux[10][44] , 
        \ADDER_IN_from_mux[10][43] , \ADDER_IN_from_mux[10][42] , 
        \ADDER_IN_from_mux[10][41] , \ADDER_IN_from_mux[10][40] , 
        \ADDER_IN_from_mux[10][39] , \ADDER_IN_from_mux[10][38] , 
        \ADDER_IN_from_mux[10][37] , \ADDER_IN_from_mux[10][36] , 
        \ADDER_IN_from_mux[10][35] , \ADDER_IN_from_mux[10][34] , 
        \ADDER_IN_from_mux[10][33] , \ADDER_IN_from_mux[10][32] , 
        \ADDER_IN_from_mux[10][31] , \ADDER_IN_from_mux[10][30] , 
        \ADDER_IN_from_mux[10][29] , \ADDER_IN_from_mux[10][28] , 
        \ADDER_IN_from_mux[10][27] , \ADDER_IN_from_mux[10][26] , 
        \ADDER_IN_from_mux[10][25] , \ADDER_IN_from_mux[10][24] , 
        \ADDER_IN_from_mux[10][23] , \ADDER_IN_from_mux[10][22] , 
        \ADDER_IN_from_mux[10][21] , \ADDER_IN_from_mux[10][20] , 
        \ADDER_IN_from_mux[10][19] , \ADDER_IN_from_mux[10][18] , 
        \ADDER_IN_from_mux[10][17] , \ADDER_IN_from_mux[10][16] , 
        \ADDER_IN_from_mux[10][15] , \ADDER_IN_from_mux[10][14] , 
        \ADDER_IN_from_mux[10][13] , \ADDER_IN_from_mux[10][12] , 
        \ADDER_IN_from_mux[10][11] , \ADDER_IN_from_mux[10][10] , 
        \ADDER_IN_from_mux[10][9] , \ADDER_IN_from_mux[10][8] , 
        \ADDER_IN_from_mux[10][7] , \ADDER_IN_from_mux[10][6] , 
        \ADDER_IN_from_mux[10][5] , \ADDER_IN_from_mux[10][4] , 
        \ADDER_IN_from_mux[10][3] , \ADDER_IN_from_mux[10][2] , 
        \ADDER_IN_from_mux[10][1] , \ADDER_IN_from_mux[10][0] }) );
  MUX81_GENERIC_NBIT64_5 MUX81_N_11 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n662, 
        n662, n662, n662, n662, n662, n662, n662, n662, n662, n662, n627, n624, 
        n618, n616, n612, n610, n606, n600, n597, n594, n588, n582, n576, n572, 
        n566, n563, n557, n554, n550, n547, n542, n538, n534, n532, n530, n527, 
        n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n672, n672, n672, n672, n673, n671, n671, n671, 
        n671, n671, n628, n625, n619, n616, n613, n610, n606, n601, n598, n594, 
        n588, n583, n576, n572, n567, n564, n557, n554, n551, n548, n542, n538, 
        n534, n531, n530, n528, n506, n521, n517, n515, n507, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[22][63] , \negative_inputs[22][62] , 
        \negative_inputs[22][61] , \negative_inputs[22][60] , 
        \negative_inputs[22][59] , \negative_inputs[22][58] , 
        \negative_inputs[22][57] , \negative_inputs[22][56] , 
        \negative_inputs[22][55] , \negative_inputs[22][54] , 
        \negative_inputs[22][53] , \negative_inputs[22][52] , 
        \negative_inputs[22][51] , \negative_inputs[22][50] , 
        \negative_inputs[22][49] , \negative_inputs[22][48] , 
        \negative_inputs[22][47] , \negative_inputs[22][46] , 
        \negative_inputs[22][45] , \negative_inputs[22][44] , 
        \negative_inputs[22][43] , \negative_inputs[22][42] , 
        \negative_inputs[22][41] , \negative_inputs[22][40] , 
        \negative_inputs[22][39] , \negative_inputs[22][38] , 
        \negative_inputs[22][37] , \negative_inputs[22][36] , 
        \negative_inputs[22][35] , \negative_inputs[22][34] , 
        \negative_inputs[22][33] , \negative_inputs[22][32] , 
        \negative_inputs[22][31] , \negative_inputs[22][30] , 
        \negative_inputs[22][29] , \negative_inputs[22][28] , 
        \negative_inputs[22][27] , \negative_inputs[22][26] , 
        \negative_inputs[22][25] , \negative_inputs[22][24] , 
        \negative_inputs[22][23] , \negative_inputs[22][22] , 
        \negative_inputs[22][21] , \negative_inputs[22][20] , 
        \negative_inputs[22][19] , \negative_inputs[22][18] , 
        \negative_inputs[22][17] , \negative_inputs[22][16] , 
        \negative_inputs[22][15] , \negative_inputs[22][14] , 
        \negative_inputs[22][13] , \negative_inputs[22][12] , 
        \negative_inputs[22][11] , \negative_inputs[22][10] , 
        \negative_inputs[22][9] , \negative_inputs[22][8] , 
        \negative_inputs[22][7] , \negative_inputs[22][6] , 
        \negative_inputs[22][5] , \negative_inputs[22][4] , 
        \negative_inputs[22][3] , \negative_inputs[22][2] , 
        \negative_inputs[22][1] , \negative_inputs[22][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[23][63] , \negative_inputs[23][62] , 
        \negative_inputs[23][61] , \negative_inputs[23][60] , 
        \negative_inputs[23][59] , \negative_inputs[23][58] , 
        \negative_inputs[23][57] , \negative_inputs[23][56] , 
        \negative_inputs[23][55] , \negative_inputs[23][54] , 
        \negative_inputs[23][53] , \negative_inputs[23][52] , 
        \negative_inputs[23][51] , \negative_inputs[23][50] , 
        \negative_inputs[23][49] , \negative_inputs[23][48] , 
        \negative_inputs[23][47] , \negative_inputs[23][46] , 
        \negative_inputs[23][45] , \negative_inputs[23][44] , 
        \negative_inputs[23][43] , \negative_inputs[23][42] , 
        \negative_inputs[23][41] , \negative_inputs[23][40] , 
        \negative_inputs[23][39] , \negative_inputs[23][38] , 
        \negative_inputs[23][37] , \negative_inputs[23][36] , 
        \negative_inputs[23][35] , \negative_inputs[23][34] , 
        \negative_inputs[23][33] , \negative_inputs[23][32] , 
        \negative_inputs[23][31] , \negative_inputs[23][30] , 
        \negative_inputs[23][29] , \negative_inputs[23][28] , 
        \negative_inputs[23][27] , \negative_inputs[23][26] , 
        \negative_inputs[23][25] , \negative_inputs[23][24] , 
        \negative_inputs[23][23] , \negative_inputs[23][22] , 
        \negative_inputs[23][21] , \negative_inputs[23][20] , 
        \negative_inputs[23][19] , \negative_inputs[23][18] , 
        \negative_inputs[23][17] , \negative_inputs[23][16] , 
        \negative_inputs[23][15] , \negative_inputs[23][14] , 
        \negative_inputs[23][13] , \negative_inputs[23][12] , 
        \negative_inputs[23][11] , \negative_inputs[23][10] , 
        \negative_inputs[23][9] , \negative_inputs[23][8] , 
        \negative_inputs[23][7] , \negative_inputs[23][6] , 
        \negative_inputs[23][5] , \negative_inputs[23][4] , 
        \negative_inputs[23][3] , \negative_inputs[23][2] , 
        \negative_inputs[23][1] , \negative_inputs[23][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[35:33]), .Y({
        \ADDER_IN_from_mux[11][63] , \ADDER_IN_from_mux[11][62] , 
        \ADDER_IN_from_mux[11][61] , \ADDER_IN_from_mux[11][60] , 
        \ADDER_IN_from_mux[11][59] , \ADDER_IN_from_mux[11][58] , 
        \ADDER_IN_from_mux[11][57] , \ADDER_IN_from_mux[11][56] , 
        \ADDER_IN_from_mux[11][55] , \ADDER_IN_from_mux[11][54] , 
        \ADDER_IN_from_mux[11][53] , \ADDER_IN_from_mux[11][52] , 
        \ADDER_IN_from_mux[11][51] , \ADDER_IN_from_mux[11][50] , 
        \ADDER_IN_from_mux[11][49] , \ADDER_IN_from_mux[11][48] , 
        \ADDER_IN_from_mux[11][47] , \ADDER_IN_from_mux[11][46] , 
        \ADDER_IN_from_mux[11][45] , \ADDER_IN_from_mux[11][44] , 
        \ADDER_IN_from_mux[11][43] , \ADDER_IN_from_mux[11][42] , 
        \ADDER_IN_from_mux[11][41] , \ADDER_IN_from_mux[11][40] , 
        \ADDER_IN_from_mux[11][39] , \ADDER_IN_from_mux[11][38] , 
        \ADDER_IN_from_mux[11][37] , \ADDER_IN_from_mux[11][36] , 
        \ADDER_IN_from_mux[11][35] , \ADDER_IN_from_mux[11][34] , 
        \ADDER_IN_from_mux[11][33] , \ADDER_IN_from_mux[11][32] , 
        \ADDER_IN_from_mux[11][31] , \ADDER_IN_from_mux[11][30] , 
        \ADDER_IN_from_mux[11][29] , \ADDER_IN_from_mux[11][28] , 
        \ADDER_IN_from_mux[11][27] , \ADDER_IN_from_mux[11][26] , 
        \ADDER_IN_from_mux[11][25] , \ADDER_IN_from_mux[11][24] , 
        \ADDER_IN_from_mux[11][23] , \ADDER_IN_from_mux[11][22] , 
        \ADDER_IN_from_mux[11][21] , \ADDER_IN_from_mux[11][20] , 
        \ADDER_IN_from_mux[11][19] , \ADDER_IN_from_mux[11][18] , 
        \ADDER_IN_from_mux[11][17] , \ADDER_IN_from_mux[11][16] , 
        \ADDER_IN_from_mux[11][15] , \ADDER_IN_from_mux[11][14] , 
        \ADDER_IN_from_mux[11][13] , \ADDER_IN_from_mux[11][12] , 
        \ADDER_IN_from_mux[11][11] , \ADDER_IN_from_mux[11][10] , 
        \ADDER_IN_from_mux[11][9] , \ADDER_IN_from_mux[11][8] , 
        \ADDER_IN_from_mux[11][7] , \ADDER_IN_from_mux[11][6] , 
        \ADDER_IN_from_mux[11][5] , \ADDER_IN_from_mux[11][4] , 
        \ADDER_IN_from_mux[11][3] , \ADDER_IN_from_mux[11][2] , 
        \ADDER_IN_from_mux[11][1] , \ADDER_IN_from_mux[11][0] }) );
  MUX81_GENERIC_NBIT64_4 MUX81_N_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n662, 
        n662, n662, n662, n662, n662, n662, n662, n662, n627, n624, n618, n616, 
        n612, n610, n606, n601, n598, n594, n588, n582, n576, n572, n567, n563, 
        n557, n553, n550, n547, n542, n538, n534, n531, n491, n527, n506, n521, 
        n517, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n671, n671, n671, n672, n671, n671, n671, n671, 
        n628, n625, n619, n616, n613, n610, n607, n601, n598, n594, n588, n583, 
        n576, n572, n567, n564, n557, n554, n551, n548, n542, n538, n534, n531, 
        n530, n528, n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[24][63] , \negative_inputs[24][62] , 
        \negative_inputs[24][61] , \negative_inputs[24][60] , 
        \negative_inputs[24][59] , \negative_inputs[24][58] , 
        \negative_inputs[24][57] , \negative_inputs[24][56] , 
        \negative_inputs[24][55] , \negative_inputs[24][54] , 
        \negative_inputs[24][53] , \negative_inputs[24][52] , 
        \negative_inputs[24][51] , \negative_inputs[24][50] , 
        \negative_inputs[24][49] , \negative_inputs[24][48] , 
        \negative_inputs[24][47] , \negative_inputs[24][46] , 
        \negative_inputs[24][45] , \negative_inputs[24][44] , 
        \negative_inputs[24][43] , \negative_inputs[24][42] , 
        \negative_inputs[24][41] , \negative_inputs[24][40] , 
        \negative_inputs[24][39] , \negative_inputs[24][38] , 
        \negative_inputs[24][37] , \negative_inputs[24][36] , 
        \negative_inputs[24][35] , \negative_inputs[24][34] , 
        \negative_inputs[24][33] , \negative_inputs[24][32] , 
        \negative_inputs[24][31] , \negative_inputs[24][30] , 
        \negative_inputs[24][29] , \negative_inputs[24][28] , 
        \negative_inputs[24][27] , \negative_inputs[24][26] , 
        \negative_inputs[24][25] , \negative_inputs[24][24] , 
        \negative_inputs[24][23] , \negative_inputs[24][22] , 
        \negative_inputs[24][21] , \negative_inputs[24][20] , 
        \negative_inputs[24][19] , \negative_inputs[24][18] , 
        \negative_inputs[24][17] , \negative_inputs[24][16] , 
        \negative_inputs[24][15] , \negative_inputs[24][14] , 
        \negative_inputs[24][13] , \negative_inputs[24][12] , 
        \negative_inputs[24][11] , \negative_inputs[24][10] , 
        \negative_inputs[24][9] , \negative_inputs[24][8] , 
        \negative_inputs[24][7] , \negative_inputs[24][6] , 
        \negative_inputs[24][5] , \negative_inputs[24][4] , 
        \negative_inputs[24][3] , \negative_inputs[24][2] , 
        \negative_inputs[24][1] , \negative_inputs[24][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[25][63] , \negative_inputs[25][62] , 
        \negative_inputs[25][61] , \negative_inputs[25][60] , 
        \negative_inputs[25][59] , \negative_inputs[25][58] , 
        \negative_inputs[25][57] , \negative_inputs[25][56] , 
        \negative_inputs[25][55] , \negative_inputs[25][54] , 
        \negative_inputs[25][53] , \negative_inputs[25][52] , 
        \negative_inputs[25][51] , \negative_inputs[25][50] , 
        \negative_inputs[25][49] , \negative_inputs[25][48] , 
        \negative_inputs[25][47] , \negative_inputs[25][46] , 
        \negative_inputs[25][45] , \negative_inputs[25][44] , 
        \negative_inputs[25][43] , \negative_inputs[25][42] , 
        \negative_inputs[25][41] , \negative_inputs[25][40] , 
        \negative_inputs[25][39] , \negative_inputs[25][38] , 
        \negative_inputs[25][37] , \negative_inputs[25][36] , 
        \negative_inputs[25][35] , \negative_inputs[25][34] , 
        \negative_inputs[25][33] , \negative_inputs[25][32] , 
        \negative_inputs[25][31] , \negative_inputs[25][30] , 
        \negative_inputs[25][29] , \negative_inputs[25][28] , 
        \negative_inputs[25][27] , \negative_inputs[25][26] , 
        \negative_inputs[25][25] , \negative_inputs[25][24] , 
        \negative_inputs[25][23] , \negative_inputs[25][22] , 
        \negative_inputs[25][21] , \negative_inputs[25][20] , 
        \negative_inputs[25][19] , \negative_inputs[25][18] , 
        \negative_inputs[25][17] , \negative_inputs[25][16] , 
        \negative_inputs[25][15] , \negative_inputs[25][14] , 
        \negative_inputs[25][13] , \negative_inputs[25][12] , 
        \negative_inputs[25][11] , \negative_inputs[25][10] , 
        \negative_inputs[25][9] , \negative_inputs[25][8] , 
        \negative_inputs[25][7] , \negative_inputs[25][6] , 
        \negative_inputs[25][5] , \negative_inputs[25][4] , 
        \negative_inputs[25][3] , \negative_inputs[25][2] , 
        \negative_inputs[25][1] , \negative_inputs[25][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[38:36]), .Y({
        \ADDER_IN_from_mux[12][63] , \ADDER_IN_from_mux[12][62] , 
        \ADDER_IN_from_mux[12][61] , \ADDER_IN_from_mux[12][60] , 
        \ADDER_IN_from_mux[12][59] , \ADDER_IN_from_mux[12][58] , 
        \ADDER_IN_from_mux[12][57] , \ADDER_IN_from_mux[12][56] , 
        \ADDER_IN_from_mux[12][55] , \ADDER_IN_from_mux[12][54] , 
        \ADDER_IN_from_mux[12][53] , \ADDER_IN_from_mux[12][52] , 
        \ADDER_IN_from_mux[12][51] , \ADDER_IN_from_mux[12][50] , 
        \ADDER_IN_from_mux[12][49] , \ADDER_IN_from_mux[12][48] , 
        \ADDER_IN_from_mux[12][47] , \ADDER_IN_from_mux[12][46] , 
        \ADDER_IN_from_mux[12][45] , \ADDER_IN_from_mux[12][44] , 
        \ADDER_IN_from_mux[12][43] , \ADDER_IN_from_mux[12][42] , 
        \ADDER_IN_from_mux[12][41] , \ADDER_IN_from_mux[12][40] , 
        \ADDER_IN_from_mux[12][39] , \ADDER_IN_from_mux[12][38] , 
        \ADDER_IN_from_mux[12][37] , \ADDER_IN_from_mux[12][36] , 
        \ADDER_IN_from_mux[12][35] , \ADDER_IN_from_mux[12][34] , 
        \ADDER_IN_from_mux[12][33] , \ADDER_IN_from_mux[12][32] , 
        \ADDER_IN_from_mux[12][31] , \ADDER_IN_from_mux[12][30] , 
        \ADDER_IN_from_mux[12][29] , \ADDER_IN_from_mux[12][28] , 
        \ADDER_IN_from_mux[12][27] , \ADDER_IN_from_mux[12][26] , 
        \ADDER_IN_from_mux[12][25] , \ADDER_IN_from_mux[12][24] , 
        \ADDER_IN_from_mux[12][23] , \ADDER_IN_from_mux[12][22] , 
        \ADDER_IN_from_mux[12][21] , \ADDER_IN_from_mux[12][20] , 
        \ADDER_IN_from_mux[12][19] , \ADDER_IN_from_mux[12][18] , 
        \ADDER_IN_from_mux[12][17] , \ADDER_IN_from_mux[12][16] , 
        \ADDER_IN_from_mux[12][15] , \ADDER_IN_from_mux[12][14] , 
        \ADDER_IN_from_mux[12][13] , \ADDER_IN_from_mux[12][12] , 
        \ADDER_IN_from_mux[12][11] , \ADDER_IN_from_mux[12][10] , 
        \ADDER_IN_from_mux[12][9] , \ADDER_IN_from_mux[12][8] , 
        \ADDER_IN_from_mux[12][7] , \ADDER_IN_from_mux[12][6] , 
        \ADDER_IN_from_mux[12][5] , \ADDER_IN_from_mux[12][4] , 
        \ADDER_IN_from_mux[12][3] , \ADDER_IN_from_mux[12][2] , 
        \ADDER_IN_from_mux[12][1] , \ADDER_IN_from_mux[12][0] }) );
  MUX81_GENERIC_NBIT64_3 MUX81_N_13 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n662, 
        n662, n662, n662, n663, n663, n663, n627, n624, n618, n616, n612, n610, 
        n606, n601, n598, n594, n588, n582, n576, n572, n567, n563, n557, n553, 
        n551, n547, n542, n538, n534, n531, n530, n527, n506, n521, n517, n515, 
        n493, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n671, n671, n670, n670, n670, n670, n628, n625, 
        n619, n616, n613, n610, n607, n601, n598, n594, n588, n583, n576, n572, 
        n567, n564, n557, n554, n551, n548, n542, n538, n535, n532, n491, n528, 
        n506, n521, n518, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[26][63] , \negative_inputs[26][62] , 
        \negative_inputs[26][61] , \negative_inputs[26][60] , 
        \negative_inputs[26][59] , \negative_inputs[26][58] , 
        \negative_inputs[26][57] , \negative_inputs[26][56] , 
        \negative_inputs[26][55] , \negative_inputs[26][54] , 
        \negative_inputs[26][53] , \negative_inputs[26][52] , 
        \negative_inputs[26][51] , \negative_inputs[26][50] , 
        \negative_inputs[26][49] , \negative_inputs[26][48] , 
        \negative_inputs[26][47] , \negative_inputs[26][46] , 
        \negative_inputs[26][45] , \negative_inputs[26][44] , 
        \negative_inputs[26][43] , \negative_inputs[26][42] , 
        \negative_inputs[26][41] , \negative_inputs[26][40] , 
        \negative_inputs[26][39] , \negative_inputs[26][38] , 
        \negative_inputs[26][37] , \negative_inputs[26][36] , 
        \negative_inputs[26][35] , \negative_inputs[26][34] , 
        \negative_inputs[26][33] , \negative_inputs[26][32] , 
        \negative_inputs[26][31] , \negative_inputs[26][30] , 
        \negative_inputs[26][29] , \negative_inputs[26][28] , 
        \negative_inputs[26][27] , \negative_inputs[26][26] , 
        \negative_inputs[26][25] , \negative_inputs[26][24] , 
        \negative_inputs[26][23] , \negative_inputs[26][22] , 
        \negative_inputs[26][21] , \negative_inputs[26][20] , 
        \negative_inputs[26][19] , \negative_inputs[26][18] , 
        \negative_inputs[26][17] , \negative_inputs[26][16] , 
        \negative_inputs[26][15] , \negative_inputs[26][14] , 
        \negative_inputs[26][13] , \negative_inputs[26][12] , 
        \negative_inputs[26][11] , \negative_inputs[26][10] , 
        \negative_inputs[26][9] , \negative_inputs[26][8] , 
        \negative_inputs[26][7] , \negative_inputs[26][6] , 
        \negative_inputs[26][5] , \negative_inputs[26][4] , 
        \negative_inputs[26][3] , \negative_inputs[26][2] , 
        \negative_inputs[26][1] , \negative_inputs[26][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[27][63] , \negative_inputs[27][62] , 
        \negative_inputs[27][61] , \negative_inputs[27][60] , 
        \negative_inputs[27][59] , \negative_inputs[27][58] , 
        \negative_inputs[27][57] , \negative_inputs[27][56] , 
        \negative_inputs[27][55] , \negative_inputs[27][54] , 
        \negative_inputs[27][53] , \negative_inputs[27][52] , 
        \negative_inputs[27][51] , \negative_inputs[27][50] , 
        \negative_inputs[27][49] , \negative_inputs[27][48] , 
        \negative_inputs[27][47] , \negative_inputs[27][46] , 
        \negative_inputs[27][45] , \negative_inputs[27][44] , 
        \negative_inputs[27][43] , \negative_inputs[27][42] , 
        \negative_inputs[27][41] , \negative_inputs[27][40] , 
        \negative_inputs[27][39] , \negative_inputs[27][38] , 
        \negative_inputs[27][37] , \negative_inputs[27][36] , 
        \negative_inputs[27][35] , \negative_inputs[27][34] , 
        \negative_inputs[27][33] , \negative_inputs[27][32] , 
        \negative_inputs[27][31] , \negative_inputs[27][30] , 
        \negative_inputs[27][29] , \negative_inputs[27][28] , 
        \negative_inputs[27][27] , \negative_inputs[27][26] , 
        \negative_inputs[27][25] , \negative_inputs[27][24] , 
        \negative_inputs[27][23] , \negative_inputs[27][22] , 
        \negative_inputs[27][21] , \negative_inputs[27][20] , 
        \negative_inputs[27][19] , \negative_inputs[27][18] , 
        \negative_inputs[27][17] , \negative_inputs[27][16] , 
        \negative_inputs[27][15] , \negative_inputs[27][14] , 
        \negative_inputs[27][13] , \negative_inputs[27][12] , 
        \negative_inputs[27][11] , \negative_inputs[27][10] , 
        \negative_inputs[27][9] , \negative_inputs[27][8] , 
        \negative_inputs[27][7] , \negative_inputs[27][6] , 
        \negative_inputs[27][5] , \negative_inputs[27][4] , 
        \negative_inputs[27][3] , \negative_inputs[27][2] , 
        \negative_inputs[27][1] , \negative_inputs[27][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[41:39]), .Y({
        \ADDER_IN_from_mux[13][63] , \ADDER_IN_from_mux[13][62] , 
        \ADDER_IN_from_mux[13][61] , \ADDER_IN_from_mux[13][60] , 
        \ADDER_IN_from_mux[13][59] , \ADDER_IN_from_mux[13][58] , 
        \ADDER_IN_from_mux[13][57] , \ADDER_IN_from_mux[13][56] , 
        \ADDER_IN_from_mux[13][55] , \ADDER_IN_from_mux[13][54] , 
        \ADDER_IN_from_mux[13][53] , \ADDER_IN_from_mux[13][52] , 
        \ADDER_IN_from_mux[13][51] , \ADDER_IN_from_mux[13][50] , 
        \ADDER_IN_from_mux[13][49] , \ADDER_IN_from_mux[13][48] , 
        \ADDER_IN_from_mux[13][47] , \ADDER_IN_from_mux[13][46] , 
        \ADDER_IN_from_mux[13][45] , \ADDER_IN_from_mux[13][44] , 
        \ADDER_IN_from_mux[13][43] , \ADDER_IN_from_mux[13][42] , 
        \ADDER_IN_from_mux[13][41] , \ADDER_IN_from_mux[13][40] , 
        \ADDER_IN_from_mux[13][39] , \ADDER_IN_from_mux[13][38] , 
        \ADDER_IN_from_mux[13][37] , \ADDER_IN_from_mux[13][36] , 
        \ADDER_IN_from_mux[13][35] , \ADDER_IN_from_mux[13][34] , 
        \ADDER_IN_from_mux[13][33] , \ADDER_IN_from_mux[13][32] , 
        \ADDER_IN_from_mux[13][31] , \ADDER_IN_from_mux[13][30] , 
        \ADDER_IN_from_mux[13][29] , \ADDER_IN_from_mux[13][28] , 
        \ADDER_IN_from_mux[13][27] , \ADDER_IN_from_mux[13][26] , 
        \ADDER_IN_from_mux[13][25] , \ADDER_IN_from_mux[13][24] , 
        \ADDER_IN_from_mux[13][23] , \ADDER_IN_from_mux[13][22] , 
        \ADDER_IN_from_mux[13][21] , \ADDER_IN_from_mux[13][20] , 
        \ADDER_IN_from_mux[13][19] , \ADDER_IN_from_mux[13][18] , 
        \ADDER_IN_from_mux[13][17] , \ADDER_IN_from_mux[13][16] , 
        \ADDER_IN_from_mux[13][15] , \ADDER_IN_from_mux[13][14] , 
        \ADDER_IN_from_mux[13][13] , \ADDER_IN_from_mux[13][12] , 
        \ADDER_IN_from_mux[13][11] , \ADDER_IN_from_mux[13][10] , 
        \ADDER_IN_from_mux[13][9] , \ADDER_IN_from_mux[13][8] , 
        \ADDER_IN_from_mux[13][7] , \ADDER_IN_from_mux[13][6] , 
        \ADDER_IN_from_mux[13][5] , \ADDER_IN_from_mux[13][4] , 
        \ADDER_IN_from_mux[13][3] , \ADDER_IN_from_mux[13][2] , 
        \ADDER_IN_from_mux[13][1] , \ADDER_IN_from_mux[13][0] }) );
  MUX81_GENERIC_NBIT64_2 MUX81_N_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n663, 
        n663, n663, n663, n663, n627, n624, n619, n616, n612, n610, n606, n601, 
        n597, n594, n588, n582, n576, n572, n566, n563, n557, n554, n551, n547, 
        n542, n537, n534, n531, n530, n527, n506, n521, n517, n515, n493, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n670, n670, n670, n670, n628, n625, n619, n616, 
        n613, n610, n607, n601, n598, n594, n588, n583, n576, n572, n567, n564, 
        n557, n554, n551, n548, n542, n538, n534, n531, n491, n528, n506, n500, 
        n518, n515, n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[28][63] , \negative_inputs[28][62] , 
        \negative_inputs[28][61] , \negative_inputs[28][60] , 
        \negative_inputs[28][59] , \negative_inputs[28][58] , 
        \negative_inputs[28][57] , \negative_inputs[28][56] , 
        \negative_inputs[28][55] , \negative_inputs[28][54] , 
        \negative_inputs[28][53] , \negative_inputs[28][52] , 
        \negative_inputs[28][51] , \negative_inputs[28][50] , 
        \negative_inputs[28][49] , \negative_inputs[28][48] , 
        \negative_inputs[28][47] , \negative_inputs[28][46] , 
        \negative_inputs[28][45] , \negative_inputs[28][44] , 
        \negative_inputs[28][43] , \negative_inputs[28][42] , 
        \negative_inputs[28][41] , \negative_inputs[28][40] , 
        \negative_inputs[28][39] , \negative_inputs[28][38] , 
        \negative_inputs[28][37] , \negative_inputs[28][36] , 
        \negative_inputs[28][35] , \negative_inputs[28][34] , 
        \negative_inputs[28][33] , \negative_inputs[28][32] , 
        \negative_inputs[28][31] , \negative_inputs[28][30] , 
        \negative_inputs[28][29] , \negative_inputs[28][28] , 
        \negative_inputs[28][27] , \negative_inputs[28][26] , 
        \negative_inputs[28][25] , \negative_inputs[28][24] , 
        \negative_inputs[28][23] , \negative_inputs[28][22] , 
        \negative_inputs[28][21] , \negative_inputs[28][20] , 
        \negative_inputs[28][19] , \negative_inputs[28][18] , 
        \negative_inputs[28][17] , \negative_inputs[28][16] , 
        \negative_inputs[28][15] , \negative_inputs[28][14] , 
        \negative_inputs[28][13] , \negative_inputs[28][12] , 
        \negative_inputs[28][11] , \negative_inputs[28][10] , 
        \negative_inputs[28][9] , \negative_inputs[28][8] , 
        \negative_inputs[28][7] , \negative_inputs[28][6] , 
        \negative_inputs[28][5] , \negative_inputs[28][4] , 
        \negative_inputs[28][3] , \negative_inputs[28][2] , 
        \negative_inputs[28][1] , \negative_inputs[28][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[29][63] , \negative_inputs[29][62] , 
        \negative_inputs[29][61] , \negative_inputs[29][60] , 
        \negative_inputs[29][59] , \negative_inputs[29][58] , 
        \negative_inputs[29][57] , \negative_inputs[29][56] , 
        \negative_inputs[29][55] , \negative_inputs[29][54] , 
        \negative_inputs[29][53] , \negative_inputs[29][52] , 
        \negative_inputs[29][51] , \negative_inputs[29][50] , 
        \negative_inputs[29][49] , \negative_inputs[29][48] , 
        \negative_inputs[29][47] , \negative_inputs[29][46] , 
        \negative_inputs[29][45] , \negative_inputs[29][44] , 
        \negative_inputs[29][43] , \negative_inputs[29][42] , 
        \negative_inputs[29][41] , \negative_inputs[29][40] , 
        \negative_inputs[29][39] , \negative_inputs[29][38] , 
        \negative_inputs[29][37] , \negative_inputs[29][36] , 
        \negative_inputs[29][35] , \negative_inputs[29][34] , 
        \negative_inputs[29][33] , \negative_inputs[29][32] , 
        \negative_inputs[29][31] , \negative_inputs[29][30] , 
        \negative_inputs[29][29] , \negative_inputs[29][28] , 
        \negative_inputs[29][27] , \negative_inputs[29][26] , 
        \negative_inputs[29][25] , \negative_inputs[29][24] , 
        \negative_inputs[29][23] , \negative_inputs[29][22] , 
        \negative_inputs[29][21] , \negative_inputs[29][20] , 
        \negative_inputs[29][19] , \negative_inputs[29][18] , 
        \negative_inputs[29][17] , \negative_inputs[29][16] , 
        \negative_inputs[29][15] , \negative_inputs[29][14] , 
        \negative_inputs[29][13] , \negative_inputs[29][12] , 
        \negative_inputs[29][11] , \negative_inputs[29][10] , 
        \negative_inputs[29][9] , \negative_inputs[29][8] , 
        \negative_inputs[29][7] , \negative_inputs[29][6] , 
        \negative_inputs[29][5] , \negative_inputs[29][4] , 
        \negative_inputs[29][3] , \negative_inputs[29][2] , 
        \negative_inputs[29][1] , \negative_inputs[29][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[44:42]), .Y({
        \ADDER_IN_from_mux[14][63] , \ADDER_IN_from_mux[14][62] , 
        \ADDER_IN_from_mux[14][61] , \ADDER_IN_from_mux[14][60] , 
        \ADDER_IN_from_mux[14][59] , \ADDER_IN_from_mux[14][58] , 
        \ADDER_IN_from_mux[14][57] , \ADDER_IN_from_mux[14][56] , 
        \ADDER_IN_from_mux[14][55] , \ADDER_IN_from_mux[14][54] , 
        \ADDER_IN_from_mux[14][53] , \ADDER_IN_from_mux[14][52] , 
        \ADDER_IN_from_mux[14][51] , \ADDER_IN_from_mux[14][50] , 
        \ADDER_IN_from_mux[14][49] , \ADDER_IN_from_mux[14][48] , 
        \ADDER_IN_from_mux[14][47] , \ADDER_IN_from_mux[14][46] , 
        \ADDER_IN_from_mux[14][45] , \ADDER_IN_from_mux[14][44] , 
        \ADDER_IN_from_mux[14][43] , \ADDER_IN_from_mux[14][42] , 
        \ADDER_IN_from_mux[14][41] , \ADDER_IN_from_mux[14][40] , 
        \ADDER_IN_from_mux[14][39] , \ADDER_IN_from_mux[14][38] , 
        \ADDER_IN_from_mux[14][37] , \ADDER_IN_from_mux[14][36] , 
        \ADDER_IN_from_mux[14][35] , \ADDER_IN_from_mux[14][34] , 
        \ADDER_IN_from_mux[14][33] , \ADDER_IN_from_mux[14][32] , 
        \ADDER_IN_from_mux[14][31] , \ADDER_IN_from_mux[14][30] , 
        \ADDER_IN_from_mux[14][29] , \ADDER_IN_from_mux[14][28] , 
        \ADDER_IN_from_mux[14][27] , \ADDER_IN_from_mux[14][26] , 
        \ADDER_IN_from_mux[14][25] , \ADDER_IN_from_mux[14][24] , 
        \ADDER_IN_from_mux[14][23] , \ADDER_IN_from_mux[14][22] , 
        \ADDER_IN_from_mux[14][21] , \ADDER_IN_from_mux[14][20] , 
        \ADDER_IN_from_mux[14][19] , \ADDER_IN_from_mux[14][18] , 
        \ADDER_IN_from_mux[14][17] , \ADDER_IN_from_mux[14][16] , 
        \ADDER_IN_from_mux[14][15] , \ADDER_IN_from_mux[14][14] , 
        \ADDER_IN_from_mux[14][13] , \ADDER_IN_from_mux[14][12] , 
        \ADDER_IN_from_mux[14][11] , \ADDER_IN_from_mux[14][10] , 
        \ADDER_IN_from_mux[14][9] , \ADDER_IN_from_mux[14][8] , 
        \ADDER_IN_from_mux[14][7] , \ADDER_IN_from_mux[14][6] , 
        \ADDER_IN_from_mux[14][5] , \ADDER_IN_from_mux[14][4] , 
        \ADDER_IN_from_mux[14][3] , \ADDER_IN_from_mux[14][2] , 
        \ADDER_IN_from_mux[14][1] , \ADDER_IN_from_mux[14][0] }) );
  MUX81_GENERIC_NBIT64_1 MUX81_N_15 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n663, 
        n663, n657, n627, n624, n618, n616, n613, n610, n606, n601, n597, n594, 
        n588, n582, n576, n572, n567, n563, n556, n554, n550, n547, n542, n537, 
        n534, n531, n530, n527, n506, n521, n517, n515, n493, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .C({n670, n666, n628, n625, n619, n616, n613, n610, 
        n606, n601, n598, n594, n588, n583, n576, n572, n567, n564, n557, n554, 
        n551, n547, n542, n537, n534, n531, n530, n527, n506, n521, n517, n515, 
        n507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({\negative_inputs[30][63] , \negative_inputs[30][62] , 
        \negative_inputs[30][61] , \negative_inputs[30][60] , 
        \negative_inputs[30][59] , \negative_inputs[30][58] , 
        \negative_inputs[30][57] , \negative_inputs[30][56] , 
        \negative_inputs[30][55] , \negative_inputs[30][54] , 
        \negative_inputs[30][53] , \negative_inputs[30][52] , 
        \negative_inputs[30][51] , \negative_inputs[30][50] , 
        \negative_inputs[30][49] , \negative_inputs[30][48] , 
        \negative_inputs[30][47] , \negative_inputs[30][46] , 
        \negative_inputs[30][45] , \negative_inputs[30][44] , 
        \negative_inputs[30][43] , \negative_inputs[30][42] , 
        \negative_inputs[30][41] , \negative_inputs[30][40] , 
        \negative_inputs[30][39] , \negative_inputs[30][38] , 
        \negative_inputs[30][37] , \negative_inputs[30][36] , 
        \negative_inputs[30][35] , \negative_inputs[30][34] , 
        \negative_inputs[30][33] , \negative_inputs[30][32] , 
        \negative_inputs[30][31] , \negative_inputs[30][30] , 
        \negative_inputs[30][29] , \negative_inputs[30][28] , 
        \negative_inputs[30][27] , \negative_inputs[30][26] , 
        \negative_inputs[30][25] , \negative_inputs[30][24] , 
        \negative_inputs[30][23] , \negative_inputs[30][22] , 
        \negative_inputs[30][21] , \negative_inputs[30][20] , 
        \negative_inputs[30][19] , \negative_inputs[30][18] , 
        \negative_inputs[30][17] , \negative_inputs[30][16] , 
        \negative_inputs[30][15] , \negative_inputs[30][14] , 
        \negative_inputs[30][13] , \negative_inputs[30][12] , 
        \negative_inputs[30][11] , \negative_inputs[30][10] , 
        \negative_inputs[30][9] , \negative_inputs[30][8] , 
        \negative_inputs[30][7] , \negative_inputs[30][6] , 
        \negative_inputs[30][5] , \negative_inputs[30][4] , 
        \negative_inputs[30][3] , \negative_inputs[30][2] , 
        \negative_inputs[30][1] , \negative_inputs[30][0] }), .F({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .G({\negative_inputs[31][63] , \negative_inputs[31][62] , 
        \negative_inputs[31][61] , \negative_inputs[31][60] , 
        \negative_inputs[31][59] , \negative_inputs[31][58] , 
        \negative_inputs[31][57] , \negative_inputs[31][56] , 
        \negative_inputs[31][55] , \negative_inputs[31][54] , 
        \negative_inputs[31][53] , \negative_inputs[31][52] , 
        \negative_inputs[31][51] , \negative_inputs[31][50] , 
        \negative_inputs[31][49] , \negative_inputs[31][48] , 
        \negative_inputs[31][47] , \negative_inputs[31][46] , 
        \negative_inputs[31][45] , \negative_inputs[31][44] , 
        \negative_inputs[31][43] , \negative_inputs[31][42] , 
        \negative_inputs[31][41] , \negative_inputs[31][40] , 
        \negative_inputs[31][39] , \negative_inputs[31][38] , 
        \negative_inputs[31][37] , \negative_inputs[31][36] , 
        \negative_inputs[31][35] , \negative_inputs[31][34] , 
        \negative_inputs[31][33] , \negative_inputs[31][32] , 
        \negative_inputs[31][31] , \negative_inputs[31][30] , 
        \negative_inputs[31][29] , \negative_inputs[31][28] , 
        \negative_inputs[31][27] , \negative_inputs[31][26] , 
        \negative_inputs[31][25] , \negative_inputs[31][24] , 
        \negative_inputs[31][23] , \negative_inputs[31][22] , 
        \negative_inputs[31][21] , \negative_inputs[31][20] , 
        \negative_inputs[31][19] , \negative_inputs[31][18] , 
        \negative_inputs[31][17] , \negative_inputs[31][16] , 
        \negative_inputs[31][15] , \negative_inputs[31][14] , 
        \negative_inputs[31][13] , \negative_inputs[31][12] , 
        \negative_inputs[31][11] , \negative_inputs[31][10] , 
        \negative_inputs[31][9] , \negative_inputs[31][8] , 
        \negative_inputs[31][7] , \negative_inputs[31][6] , 
        \negative_inputs[31][5] , \negative_inputs[31][4] , 
        \negative_inputs[31][3] , \negative_inputs[31][2] , 
        \negative_inputs[31][1] , \negative_inputs[31][0] }), .H({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL(Encoder_out[47:45]), .Y({
        \ADDER_IN_from_mux[15][63] , \ADDER_IN_from_mux[15][62] , 
        \ADDER_IN_from_mux[15][61] , \ADDER_IN_from_mux[15][60] , 
        \ADDER_IN_from_mux[15][59] , \ADDER_IN_from_mux[15][58] , 
        \ADDER_IN_from_mux[15][57] , \ADDER_IN_from_mux[15][56] , 
        \ADDER_IN_from_mux[15][55] , \ADDER_IN_from_mux[15][54] , 
        \ADDER_IN_from_mux[15][53] , \ADDER_IN_from_mux[15][52] , 
        \ADDER_IN_from_mux[15][51] , \ADDER_IN_from_mux[15][50] , 
        \ADDER_IN_from_mux[15][49] , \ADDER_IN_from_mux[15][48] , 
        \ADDER_IN_from_mux[15][47] , \ADDER_IN_from_mux[15][46] , 
        \ADDER_IN_from_mux[15][45] , \ADDER_IN_from_mux[15][44] , 
        \ADDER_IN_from_mux[15][43] , \ADDER_IN_from_mux[15][42] , 
        \ADDER_IN_from_mux[15][41] , \ADDER_IN_from_mux[15][40] , 
        \ADDER_IN_from_mux[15][39] , \ADDER_IN_from_mux[15][38] , 
        \ADDER_IN_from_mux[15][37] , \ADDER_IN_from_mux[15][36] , 
        \ADDER_IN_from_mux[15][35] , \ADDER_IN_from_mux[15][34] , 
        \ADDER_IN_from_mux[15][33] , \ADDER_IN_from_mux[15][32] , 
        \ADDER_IN_from_mux[15][31] , \ADDER_IN_from_mux[15][30] , 
        \ADDER_IN_from_mux[15][29] , \ADDER_IN_from_mux[15][28] , 
        \ADDER_IN_from_mux[15][27] , \ADDER_IN_from_mux[15][26] , 
        \ADDER_IN_from_mux[15][25] , \ADDER_IN_from_mux[15][24] , 
        \ADDER_IN_from_mux[15][23] , \ADDER_IN_from_mux[15][22] , 
        \ADDER_IN_from_mux[15][21] , \ADDER_IN_from_mux[15][20] , 
        \ADDER_IN_from_mux[15][19] , \ADDER_IN_from_mux[15][18] , 
        \ADDER_IN_from_mux[15][17] , \ADDER_IN_from_mux[15][16] , 
        \ADDER_IN_from_mux[15][15] , \ADDER_IN_from_mux[15][14] , 
        \ADDER_IN_from_mux[15][13] , \ADDER_IN_from_mux[15][12] , 
        \ADDER_IN_from_mux[15][11] , \ADDER_IN_from_mux[15][10] , 
        \ADDER_IN_from_mux[15][9] , \ADDER_IN_from_mux[15][8] , 
        \ADDER_IN_from_mux[15][7] , \ADDER_IN_from_mux[15][6] , 
        \ADDER_IN_from_mux[15][5] , \ADDER_IN_from_mux[15][4] , 
        \ADDER_IN_from_mux[15][3] , \ADDER_IN_from_mux[15][2] , 
        \ADDER_IN_from_mux[15][1] , \ADDER_IN_from_mux[15][0] }) );
  RCA_NBIT64_0 first_adder ( .A({\ADDER_IN_from_mux[0][63] , 
        \ADDER_IN_from_mux[0][62] , \ADDER_IN_from_mux[0][61] , 
        \ADDER_IN_from_mux[0][60] , \ADDER_IN_from_mux[0][59] , 
        \ADDER_IN_from_mux[0][58] , \ADDER_IN_from_mux[0][57] , 
        \ADDER_IN_from_mux[0][56] , \ADDER_IN_from_mux[0][55] , 
        \ADDER_IN_from_mux[0][54] , \ADDER_IN_from_mux[0][53] , 
        \ADDER_IN_from_mux[0][52] , \ADDER_IN_from_mux[0][51] , 
        \ADDER_IN_from_mux[0][50] , \ADDER_IN_from_mux[0][49] , 
        \ADDER_IN_from_mux[0][48] , \ADDER_IN_from_mux[0][47] , 
        \ADDER_IN_from_mux[0][46] , \ADDER_IN_from_mux[0][45] , 
        \ADDER_IN_from_mux[0][44] , \ADDER_IN_from_mux[0][43] , 
        \ADDER_IN_from_mux[0][42] , \ADDER_IN_from_mux[0][41] , 
        \ADDER_IN_from_mux[0][40] , \ADDER_IN_from_mux[0][39] , 
        \ADDER_IN_from_mux[0][38] , \ADDER_IN_from_mux[0][37] , 
        \ADDER_IN_from_mux[0][36] , \ADDER_IN_from_mux[0][35] , 
        \ADDER_IN_from_mux[0][34] , \ADDER_IN_from_mux[0][33] , 
        \ADDER_IN_from_mux[0][32] , \ADDER_IN_from_mux[0][31] , 
        \ADDER_IN_from_mux[0][30] , \ADDER_IN_from_mux[0][29] , 
        \ADDER_IN_from_mux[0][28] , \ADDER_IN_from_mux[0][27] , 
        \ADDER_IN_from_mux[0][26] , \ADDER_IN_from_mux[0][25] , 
        \ADDER_IN_from_mux[0][24] , \ADDER_IN_from_mux[0][23] , 
        \ADDER_IN_from_mux[0][22] , \ADDER_IN_from_mux[0][21] , 
        \ADDER_IN_from_mux[0][20] , \ADDER_IN_from_mux[0][19] , 
        \ADDER_IN_from_mux[0][18] , \ADDER_IN_from_mux[0][17] , 
        \ADDER_IN_from_mux[0][16] , \ADDER_IN_from_mux[0][15] , 
        \ADDER_IN_from_mux[0][14] , \ADDER_IN_from_mux[0][13] , 
        \ADDER_IN_from_mux[0][12] , \ADDER_IN_from_mux[0][11] , 
        \ADDER_IN_from_mux[0][10] , \ADDER_IN_from_mux[0][9] , 
        \ADDER_IN_from_mux[0][8] , \ADDER_IN_from_mux[0][7] , 
        \ADDER_IN_from_mux[0][6] , \ADDER_IN_from_mux[0][5] , 
        \ADDER_IN_from_mux[0][4] , \ADDER_IN_from_mux[0][3] , 
        \ADDER_IN_from_mux[0][2] , \ADDER_IN_from_mux[0][1] , 
        \ADDER_IN_from_mux[0][0] }), .B({\ADDER_IN_from_mux[1][63] , 
        \ADDER_IN_from_mux[1][62] , \ADDER_IN_from_mux[1][61] , 
        \ADDER_IN_from_mux[1][60] , \ADDER_IN_from_mux[1][59] , 
        \ADDER_IN_from_mux[1][58] , \ADDER_IN_from_mux[1][57] , 
        \ADDER_IN_from_mux[1][56] , \ADDER_IN_from_mux[1][55] , 
        \ADDER_IN_from_mux[1][54] , \ADDER_IN_from_mux[1][53] , 
        \ADDER_IN_from_mux[1][52] , \ADDER_IN_from_mux[1][51] , 
        \ADDER_IN_from_mux[1][50] , \ADDER_IN_from_mux[1][49] , 
        \ADDER_IN_from_mux[1][48] , \ADDER_IN_from_mux[1][47] , 
        \ADDER_IN_from_mux[1][46] , \ADDER_IN_from_mux[1][45] , 
        \ADDER_IN_from_mux[1][44] , \ADDER_IN_from_mux[1][43] , 
        \ADDER_IN_from_mux[1][42] , \ADDER_IN_from_mux[1][41] , 
        \ADDER_IN_from_mux[1][40] , \ADDER_IN_from_mux[1][39] , 
        \ADDER_IN_from_mux[1][38] , \ADDER_IN_from_mux[1][37] , 
        \ADDER_IN_from_mux[1][36] , \ADDER_IN_from_mux[1][35] , 
        \ADDER_IN_from_mux[1][34] , \ADDER_IN_from_mux[1][33] , 
        \ADDER_IN_from_mux[1][32] , \ADDER_IN_from_mux[1][31] , 
        \ADDER_IN_from_mux[1][30] , \ADDER_IN_from_mux[1][29] , 
        \ADDER_IN_from_mux[1][28] , \ADDER_IN_from_mux[1][27] , 
        \ADDER_IN_from_mux[1][26] , \ADDER_IN_from_mux[1][25] , 
        \ADDER_IN_from_mux[1][24] , \ADDER_IN_from_mux[1][23] , 
        \ADDER_IN_from_mux[1][22] , \ADDER_IN_from_mux[1][21] , 
        \ADDER_IN_from_mux[1][20] , \ADDER_IN_from_mux[1][19] , 
        \ADDER_IN_from_mux[1][18] , \ADDER_IN_from_mux[1][17] , 
        \ADDER_IN_from_mux[1][16] , \ADDER_IN_from_mux[1][15] , 
        \ADDER_IN_from_mux[1][14] , \ADDER_IN_from_mux[1][13] , 
        \ADDER_IN_from_mux[1][12] , \ADDER_IN_from_mux[1][11] , 
        \ADDER_IN_from_mux[1][10] , \ADDER_IN_from_mux[1][9] , 
        \ADDER_IN_from_mux[1][8] , \ADDER_IN_from_mux[1][7] , 
        \ADDER_IN_from_mux[1][6] , \ADDER_IN_from_mux[1][5] , 
        \ADDER_IN_from_mux[1][4] , \ADDER_IN_from_mux[1][3] , 
        \ADDER_IN_from_mux[1][2] , \ADDER_IN_from_mux[1][1] , 
        \ADDER_IN_from_mux[1][0] }), .S({\ADDER_IN_from_sum[0][63] , 
        \ADDER_IN_from_sum[0][62] , \ADDER_IN_from_sum[0][61] , 
        \ADDER_IN_from_sum[0][60] , \ADDER_IN_from_sum[0][59] , 
        \ADDER_IN_from_sum[0][58] , \ADDER_IN_from_sum[0][57] , 
        \ADDER_IN_from_sum[0][56] , \ADDER_IN_from_sum[0][55] , 
        \ADDER_IN_from_sum[0][54] , \ADDER_IN_from_sum[0][53] , 
        \ADDER_IN_from_sum[0][52] , \ADDER_IN_from_sum[0][51] , 
        \ADDER_IN_from_sum[0][50] , \ADDER_IN_from_sum[0][49] , 
        \ADDER_IN_from_sum[0][48] , \ADDER_IN_from_sum[0][47] , 
        \ADDER_IN_from_sum[0][46] , \ADDER_IN_from_sum[0][45] , 
        \ADDER_IN_from_sum[0][44] , \ADDER_IN_from_sum[0][43] , 
        \ADDER_IN_from_sum[0][42] , \ADDER_IN_from_sum[0][41] , 
        \ADDER_IN_from_sum[0][40] , \ADDER_IN_from_sum[0][39] , 
        \ADDER_IN_from_sum[0][38] , \ADDER_IN_from_sum[0][37] , 
        \ADDER_IN_from_sum[0][36] , \ADDER_IN_from_sum[0][35] , 
        \ADDER_IN_from_sum[0][34] , \ADDER_IN_from_sum[0][33] , 
        \ADDER_IN_from_sum[0][32] , \ADDER_IN_from_sum[0][31] , 
        \ADDER_IN_from_sum[0][30] , \ADDER_IN_from_sum[0][29] , 
        \ADDER_IN_from_sum[0][28] , \ADDER_IN_from_sum[0][27] , 
        \ADDER_IN_from_sum[0][26] , \ADDER_IN_from_sum[0][25] , 
        \ADDER_IN_from_sum[0][24] , \ADDER_IN_from_sum[0][23] , 
        \ADDER_IN_from_sum[0][22] , \ADDER_IN_from_sum[0][21] , 
        \ADDER_IN_from_sum[0][20] , \ADDER_IN_from_sum[0][19] , 
        \ADDER_IN_from_sum[0][18] , \ADDER_IN_from_sum[0][17] , 
        \ADDER_IN_from_sum[0][16] , \ADDER_IN_from_sum[0][15] , 
        \ADDER_IN_from_sum[0][14] , \ADDER_IN_from_sum[0][13] , 
        \ADDER_IN_from_sum[0][12] , \ADDER_IN_from_sum[0][11] , 
        \ADDER_IN_from_sum[0][10] , \ADDER_IN_from_sum[0][9] , 
        \ADDER_IN_from_sum[0][8] , \ADDER_IN_from_sum[0][7] , 
        \ADDER_IN_from_sum[0][6] , \ADDER_IN_from_sum[0][5] , 
        \ADDER_IN_from_sum[0][4] , \ADDER_IN_from_sum[0][3] , 
        \ADDER_IN_from_sum[0][2] , \ADDER_IN_from_sum[0][1] , 
        \ADDER_IN_from_sum[0][0] }) );
  RCA_NBIT64_14 RCA_n_0 ( .A({\ADDER_IN_from_sum[0][63] , 
        \ADDER_IN_from_sum[0][62] , \ADDER_IN_from_sum[0][61] , 
        \ADDER_IN_from_sum[0][60] , \ADDER_IN_from_sum[0][59] , 
        \ADDER_IN_from_sum[0][58] , \ADDER_IN_from_sum[0][57] , 
        \ADDER_IN_from_sum[0][56] , \ADDER_IN_from_sum[0][55] , 
        \ADDER_IN_from_sum[0][54] , \ADDER_IN_from_sum[0][53] , 
        \ADDER_IN_from_sum[0][52] , \ADDER_IN_from_sum[0][51] , 
        \ADDER_IN_from_sum[0][50] , \ADDER_IN_from_sum[0][49] , 
        \ADDER_IN_from_sum[0][48] , \ADDER_IN_from_sum[0][47] , 
        \ADDER_IN_from_sum[0][46] , \ADDER_IN_from_sum[0][45] , 
        \ADDER_IN_from_sum[0][44] , \ADDER_IN_from_sum[0][43] , 
        \ADDER_IN_from_sum[0][42] , \ADDER_IN_from_sum[0][41] , 
        \ADDER_IN_from_sum[0][40] , \ADDER_IN_from_sum[0][39] , 
        \ADDER_IN_from_sum[0][38] , \ADDER_IN_from_sum[0][37] , 
        \ADDER_IN_from_sum[0][36] , \ADDER_IN_from_sum[0][35] , 
        \ADDER_IN_from_sum[0][34] , \ADDER_IN_from_sum[0][33] , 
        \ADDER_IN_from_sum[0][32] , \ADDER_IN_from_sum[0][31] , 
        \ADDER_IN_from_sum[0][30] , \ADDER_IN_from_sum[0][29] , 
        \ADDER_IN_from_sum[0][28] , \ADDER_IN_from_sum[0][27] , 
        \ADDER_IN_from_sum[0][26] , \ADDER_IN_from_sum[0][25] , 
        \ADDER_IN_from_sum[0][24] , \ADDER_IN_from_sum[0][23] , 
        \ADDER_IN_from_sum[0][22] , \ADDER_IN_from_sum[0][21] , 
        \ADDER_IN_from_sum[0][20] , \ADDER_IN_from_sum[0][19] , 
        \ADDER_IN_from_sum[0][18] , \ADDER_IN_from_sum[0][17] , 
        \ADDER_IN_from_sum[0][16] , \ADDER_IN_from_sum[0][15] , 
        \ADDER_IN_from_sum[0][14] , \ADDER_IN_from_sum[0][13] , 
        \ADDER_IN_from_sum[0][12] , \ADDER_IN_from_sum[0][11] , 
        \ADDER_IN_from_sum[0][10] , \ADDER_IN_from_sum[0][9] , 
        \ADDER_IN_from_sum[0][8] , \ADDER_IN_from_sum[0][7] , 
        \ADDER_IN_from_sum[0][6] , \ADDER_IN_from_sum[0][5] , 
        \ADDER_IN_from_sum[0][4] , \ADDER_IN_from_sum[0][3] , 
        \ADDER_IN_from_sum[0][2] , \ADDER_IN_from_sum[0][1] , 
        \ADDER_IN_from_sum[0][0] }), .B({\ADDER_IN_from_mux[2][63] , 
        \ADDER_IN_from_mux[2][62] , \ADDER_IN_from_mux[2][61] , 
        \ADDER_IN_from_mux[2][60] , \ADDER_IN_from_mux[2][59] , 
        \ADDER_IN_from_mux[2][58] , \ADDER_IN_from_mux[2][57] , 
        \ADDER_IN_from_mux[2][56] , \ADDER_IN_from_mux[2][55] , 
        \ADDER_IN_from_mux[2][54] , \ADDER_IN_from_mux[2][53] , 
        \ADDER_IN_from_mux[2][52] , \ADDER_IN_from_mux[2][51] , 
        \ADDER_IN_from_mux[2][50] , \ADDER_IN_from_mux[2][49] , 
        \ADDER_IN_from_mux[2][48] , \ADDER_IN_from_mux[2][47] , 
        \ADDER_IN_from_mux[2][46] , \ADDER_IN_from_mux[2][45] , 
        \ADDER_IN_from_mux[2][44] , \ADDER_IN_from_mux[2][43] , 
        \ADDER_IN_from_mux[2][42] , \ADDER_IN_from_mux[2][41] , 
        \ADDER_IN_from_mux[2][40] , \ADDER_IN_from_mux[2][39] , 
        \ADDER_IN_from_mux[2][38] , \ADDER_IN_from_mux[2][37] , 
        \ADDER_IN_from_mux[2][36] , \ADDER_IN_from_mux[2][35] , 
        \ADDER_IN_from_mux[2][34] , \ADDER_IN_from_mux[2][33] , 
        \ADDER_IN_from_mux[2][32] , \ADDER_IN_from_mux[2][31] , 
        \ADDER_IN_from_mux[2][30] , \ADDER_IN_from_mux[2][29] , 
        \ADDER_IN_from_mux[2][28] , \ADDER_IN_from_mux[2][27] , 
        \ADDER_IN_from_mux[2][26] , \ADDER_IN_from_mux[2][25] , 
        \ADDER_IN_from_mux[2][24] , \ADDER_IN_from_mux[2][23] , 
        \ADDER_IN_from_mux[2][22] , \ADDER_IN_from_mux[2][21] , 
        \ADDER_IN_from_mux[2][20] , \ADDER_IN_from_mux[2][19] , 
        \ADDER_IN_from_mux[2][18] , \ADDER_IN_from_mux[2][17] , 
        \ADDER_IN_from_mux[2][16] , \ADDER_IN_from_mux[2][15] , 
        \ADDER_IN_from_mux[2][14] , \ADDER_IN_from_mux[2][13] , 
        \ADDER_IN_from_mux[2][12] , \ADDER_IN_from_mux[2][11] , 
        \ADDER_IN_from_mux[2][10] , \ADDER_IN_from_mux[2][9] , 
        \ADDER_IN_from_mux[2][8] , \ADDER_IN_from_mux[2][7] , 
        \ADDER_IN_from_mux[2][6] , \ADDER_IN_from_mux[2][5] , 
        \ADDER_IN_from_mux[2][4] , \ADDER_IN_from_mux[2][3] , 
        \ADDER_IN_from_mux[2][2] , \ADDER_IN_from_mux[2][1] , 
        \ADDER_IN_from_mux[2][0] }), .S({\ADDER_IN_from_sum[1][63] , 
        \ADDER_IN_from_sum[1][62] , \ADDER_IN_from_sum[1][61] , 
        \ADDER_IN_from_sum[1][60] , \ADDER_IN_from_sum[1][59] , 
        \ADDER_IN_from_sum[1][58] , \ADDER_IN_from_sum[1][57] , 
        \ADDER_IN_from_sum[1][56] , \ADDER_IN_from_sum[1][55] , 
        \ADDER_IN_from_sum[1][54] , \ADDER_IN_from_sum[1][53] , 
        \ADDER_IN_from_sum[1][52] , \ADDER_IN_from_sum[1][51] , 
        \ADDER_IN_from_sum[1][50] , \ADDER_IN_from_sum[1][49] , 
        \ADDER_IN_from_sum[1][48] , \ADDER_IN_from_sum[1][47] , 
        \ADDER_IN_from_sum[1][46] , \ADDER_IN_from_sum[1][45] , 
        \ADDER_IN_from_sum[1][44] , \ADDER_IN_from_sum[1][43] , 
        \ADDER_IN_from_sum[1][42] , \ADDER_IN_from_sum[1][41] , 
        \ADDER_IN_from_sum[1][40] , \ADDER_IN_from_sum[1][39] , 
        \ADDER_IN_from_sum[1][38] , \ADDER_IN_from_sum[1][37] , 
        \ADDER_IN_from_sum[1][36] , \ADDER_IN_from_sum[1][35] , 
        \ADDER_IN_from_sum[1][34] , \ADDER_IN_from_sum[1][33] , 
        \ADDER_IN_from_sum[1][32] , \ADDER_IN_from_sum[1][31] , 
        \ADDER_IN_from_sum[1][30] , \ADDER_IN_from_sum[1][29] , 
        \ADDER_IN_from_sum[1][28] , \ADDER_IN_from_sum[1][27] , 
        \ADDER_IN_from_sum[1][26] , \ADDER_IN_from_sum[1][25] , 
        \ADDER_IN_from_sum[1][24] , \ADDER_IN_from_sum[1][23] , 
        \ADDER_IN_from_sum[1][22] , \ADDER_IN_from_sum[1][21] , 
        \ADDER_IN_from_sum[1][20] , \ADDER_IN_from_sum[1][19] , 
        \ADDER_IN_from_sum[1][18] , \ADDER_IN_from_sum[1][17] , 
        \ADDER_IN_from_sum[1][16] , \ADDER_IN_from_sum[1][15] , 
        \ADDER_IN_from_sum[1][14] , \ADDER_IN_from_sum[1][13] , 
        \ADDER_IN_from_sum[1][12] , \ADDER_IN_from_sum[1][11] , 
        \ADDER_IN_from_sum[1][10] , \ADDER_IN_from_sum[1][9] , 
        \ADDER_IN_from_sum[1][8] , \ADDER_IN_from_sum[1][7] , 
        \ADDER_IN_from_sum[1][6] , \ADDER_IN_from_sum[1][5] , 
        \ADDER_IN_from_sum[1][4] , \ADDER_IN_from_sum[1][3] , 
        \ADDER_IN_from_sum[1][2] , \ADDER_IN_from_sum[1][1] , 
        \ADDER_IN_from_sum[1][0] }) );
  RCA_NBIT64_13 RCA_n_1 ( .A({\ADDER_IN_from_sum[1][63] , 
        \ADDER_IN_from_sum[1][62] , \ADDER_IN_from_sum[1][61] , 
        \ADDER_IN_from_sum[1][60] , \ADDER_IN_from_sum[1][59] , 
        \ADDER_IN_from_sum[1][58] , \ADDER_IN_from_sum[1][57] , 
        \ADDER_IN_from_sum[1][56] , \ADDER_IN_from_sum[1][55] , 
        \ADDER_IN_from_sum[1][54] , \ADDER_IN_from_sum[1][53] , 
        \ADDER_IN_from_sum[1][52] , \ADDER_IN_from_sum[1][51] , 
        \ADDER_IN_from_sum[1][50] , \ADDER_IN_from_sum[1][49] , 
        \ADDER_IN_from_sum[1][48] , \ADDER_IN_from_sum[1][47] , 
        \ADDER_IN_from_sum[1][46] , \ADDER_IN_from_sum[1][45] , 
        \ADDER_IN_from_sum[1][44] , \ADDER_IN_from_sum[1][43] , 
        \ADDER_IN_from_sum[1][42] , \ADDER_IN_from_sum[1][41] , 
        \ADDER_IN_from_sum[1][40] , \ADDER_IN_from_sum[1][39] , 
        \ADDER_IN_from_sum[1][38] , \ADDER_IN_from_sum[1][37] , 
        \ADDER_IN_from_sum[1][36] , \ADDER_IN_from_sum[1][35] , 
        \ADDER_IN_from_sum[1][34] , \ADDER_IN_from_sum[1][33] , 
        \ADDER_IN_from_sum[1][32] , \ADDER_IN_from_sum[1][31] , 
        \ADDER_IN_from_sum[1][30] , \ADDER_IN_from_sum[1][29] , 
        \ADDER_IN_from_sum[1][28] , \ADDER_IN_from_sum[1][27] , 
        \ADDER_IN_from_sum[1][26] , \ADDER_IN_from_sum[1][25] , 
        \ADDER_IN_from_sum[1][24] , \ADDER_IN_from_sum[1][23] , 
        \ADDER_IN_from_sum[1][22] , \ADDER_IN_from_sum[1][21] , 
        \ADDER_IN_from_sum[1][20] , \ADDER_IN_from_sum[1][19] , 
        \ADDER_IN_from_sum[1][18] , \ADDER_IN_from_sum[1][17] , 
        \ADDER_IN_from_sum[1][16] , \ADDER_IN_from_sum[1][15] , 
        \ADDER_IN_from_sum[1][14] , \ADDER_IN_from_sum[1][13] , 
        \ADDER_IN_from_sum[1][12] , \ADDER_IN_from_sum[1][11] , 
        \ADDER_IN_from_sum[1][10] , \ADDER_IN_from_sum[1][9] , 
        \ADDER_IN_from_sum[1][8] , \ADDER_IN_from_sum[1][7] , 
        \ADDER_IN_from_sum[1][6] , \ADDER_IN_from_sum[1][5] , 
        \ADDER_IN_from_sum[1][4] , \ADDER_IN_from_sum[1][3] , 
        \ADDER_IN_from_sum[1][2] , \ADDER_IN_from_sum[1][1] , 
        \ADDER_IN_from_sum[1][0] }), .B({\ADDER_IN_from_mux[3][63] , 
        \ADDER_IN_from_mux[3][62] , \ADDER_IN_from_mux[3][61] , 
        \ADDER_IN_from_mux[3][60] , \ADDER_IN_from_mux[3][59] , 
        \ADDER_IN_from_mux[3][58] , \ADDER_IN_from_mux[3][57] , 
        \ADDER_IN_from_mux[3][56] , \ADDER_IN_from_mux[3][55] , 
        \ADDER_IN_from_mux[3][54] , \ADDER_IN_from_mux[3][53] , 
        \ADDER_IN_from_mux[3][52] , \ADDER_IN_from_mux[3][51] , 
        \ADDER_IN_from_mux[3][50] , \ADDER_IN_from_mux[3][49] , 
        \ADDER_IN_from_mux[3][48] , \ADDER_IN_from_mux[3][47] , 
        \ADDER_IN_from_mux[3][46] , \ADDER_IN_from_mux[3][45] , 
        \ADDER_IN_from_mux[3][44] , \ADDER_IN_from_mux[3][43] , 
        \ADDER_IN_from_mux[3][42] , \ADDER_IN_from_mux[3][41] , 
        \ADDER_IN_from_mux[3][40] , \ADDER_IN_from_mux[3][39] , 
        \ADDER_IN_from_mux[3][38] , \ADDER_IN_from_mux[3][37] , 
        \ADDER_IN_from_mux[3][36] , \ADDER_IN_from_mux[3][35] , 
        \ADDER_IN_from_mux[3][34] , \ADDER_IN_from_mux[3][33] , 
        \ADDER_IN_from_mux[3][32] , \ADDER_IN_from_mux[3][31] , 
        \ADDER_IN_from_mux[3][30] , \ADDER_IN_from_mux[3][29] , 
        \ADDER_IN_from_mux[3][28] , \ADDER_IN_from_mux[3][27] , 
        \ADDER_IN_from_mux[3][26] , \ADDER_IN_from_mux[3][25] , 
        \ADDER_IN_from_mux[3][24] , \ADDER_IN_from_mux[3][23] , 
        \ADDER_IN_from_mux[3][22] , \ADDER_IN_from_mux[3][21] , 
        \ADDER_IN_from_mux[3][20] , \ADDER_IN_from_mux[3][19] , 
        \ADDER_IN_from_mux[3][18] , \ADDER_IN_from_mux[3][17] , 
        \ADDER_IN_from_mux[3][16] , \ADDER_IN_from_mux[3][15] , 
        \ADDER_IN_from_mux[3][14] , \ADDER_IN_from_mux[3][13] , 
        \ADDER_IN_from_mux[3][12] , \ADDER_IN_from_mux[3][11] , 
        \ADDER_IN_from_mux[3][10] , \ADDER_IN_from_mux[3][9] , 
        \ADDER_IN_from_mux[3][8] , \ADDER_IN_from_mux[3][7] , 
        \ADDER_IN_from_mux[3][6] , \ADDER_IN_from_mux[3][5] , 
        \ADDER_IN_from_mux[3][4] , \ADDER_IN_from_mux[3][3] , 
        \ADDER_IN_from_mux[3][2] , \ADDER_IN_from_mux[3][1] , 
        \ADDER_IN_from_mux[3][0] }), .S({\ADDER_IN_from_sum[2][63] , 
        \ADDER_IN_from_sum[2][62] , \ADDER_IN_from_sum[2][61] , 
        \ADDER_IN_from_sum[2][60] , \ADDER_IN_from_sum[2][59] , 
        \ADDER_IN_from_sum[2][58] , \ADDER_IN_from_sum[2][57] , 
        \ADDER_IN_from_sum[2][56] , \ADDER_IN_from_sum[2][55] , 
        \ADDER_IN_from_sum[2][54] , \ADDER_IN_from_sum[2][53] , 
        \ADDER_IN_from_sum[2][52] , \ADDER_IN_from_sum[2][51] , 
        \ADDER_IN_from_sum[2][50] , \ADDER_IN_from_sum[2][49] , 
        \ADDER_IN_from_sum[2][48] , \ADDER_IN_from_sum[2][47] , 
        \ADDER_IN_from_sum[2][46] , \ADDER_IN_from_sum[2][45] , 
        \ADDER_IN_from_sum[2][44] , \ADDER_IN_from_sum[2][43] , 
        \ADDER_IN_from_sum[2][42] , \ADDER_IN_from_sum[2][41] , 
        \ADDER_IN_from_sum[2][40] , \ADDER_IN_from_sum[2][39] , 
        \ADDER_IN_from_sum[2][38] , \ADDER_IN_from_sum[2][37] , 
        \ADDER_IN_from_sum[2][36] , \ADDER_IN_from_sum[2][35] , 
        \ADDER_IN_from_sum[2][34] , \ADDER_IN_from_sum[2][33] , 
        \ADDER_IN_from_sum[2][32] , \ADDER_IN_from_sum[2][31] , 
        \ADDER_IN_from_sum[2][30] , \ADDER_IN_from_sum[2][29] , 
        \ADDER_IN_from_sum[2][28] , \ADDER_IN_from_sum[2][27] , 
        \ADDER_IN_from_sum[2][26] , \ADDER_IN_from_sum[2][25] , 
        \ADDER_IN_from_sum[2][24] , \ADDER_IN_from_sum[2][23] , 
        \ADDER_IN_from_sum[2][22] , \ADDER_IN_from_sum[2][21] , 
        \ADDER_IN_from_sum[2][20] , \ADDER_IN_from_sum[2][19] , 
        \ADDER_IN_from_sum[2][18] , \ADDER_IN_from_sum[2][17] , 
        \ADDER_IN_from_sum[2][16] , \ADDER_IN_from_sum[2][15] , 
        \ADDER_IN_from_sum[2][14] , \ADDER_IN_from_sum[2][13] , 
        \ADDER_IN_from_sum[2][12] , \ADDER_IN_from_sum[2][11] , 
        \ADDER_IN_from_sum[2][10] , \ADDER_IN_from_sum[2][9] , 
        \ADDER_IN_from_sum[2][8] , \ADDER_IN_from_sum[2][7] , 
        \ADDER_IN_from_sum[2][6] , \ADDER_IN_from_sum[2][5] , 
        \ADDER_IN_from_sum[2][4] , \ADDER_IN_from_sum[2][3] , 
        \ADDER_IN_from_sum[2][2] , \ADDER_IN_from_sum[2][1] , 
        \ADDER_IN_from_sum[2][0] }) );
  RCA_NBIT64_12 RCA_n_2 ( .A({\ADDER_IN_from_sum[2][63] , 
        \ADDER_IN_from_sum[2][62] , \ADDER_IN_from_sum[2][61] , 
        \ADDER_IN_from_sum[2][60] , \ADDER_IN_from_sum[2][59] , 
        \ADDER_IN_from_sum[2][58] , \ADDER_IN_from_sum[2][57] , 
        \ADDER_IN_from_sum[2][56] , \ADDER_IN_from_sum[2][55] , 
        \ADDER_IN_from_sum[2][54] , \ADDER_IN_from_sum[2][53] , 
        \ADDER_IN_from_sum[2][52] , \ADDER_IN_from_sum[2][51] , 
        \ADDER_IN_from_sum[2][50] , \ADDER_IN_from_sum[2][49] , 
        \ADDER_IN_from_sum[2][48] , \ADDER_IN_from_sum[2][47] , 
        \ADDER_IN_from_sum[2][46] , \ADDER_IN_from_sum[2][45] , 
        \ADDER_IN_from_sum[2][44] , \ADDER_IN_from_sum[2][43] , 
        \ADDER_IN_from_sum[2][42] , \ADDER_IN_from_sum[2][41] , 
        \ADDER_IN_from_sum[2][40] , \ADDER_IN_from_sum[2][39] , 
        \ADDER_IN_from_sum[2][38] , \ADDER_IN_from_sum[2][37] , 
        \ADDER_IN_from_sum[2][36] , \ADDER_IN_from_sum[2][35] , 
        \ADDER_IN_from_sum[2][34] , \ADDER_IN_from_sum[2][33] , 
        \ADDER_IN_from_sum[2][32] , \ADDER_IN_from_sum[2][31] , 
        \ADDER_IN_from_sum[2][30] , \ADDER_IN_from_sum[2][29] , 
        \ADDER_IN_from_sum[2][28] , \ADDER_IN_from_sum[2][27] , 
        \ADDER_IN_from_sum[2][26] , \ADDER_IN_from_sum[2][25] , 
        \ADDER_IN_from_sum[2][24] , \ADDER_IN_from_sum[2][23] , 
        \ADDER_IN_from_sum[2][22] , \ADDER_IN_from_sum[2][21] , 
        \ADDER_IN_from_sum[2][20] , \ADDER_IN_from_sum[2][19] , 
        \ADDER_IN_from_sum[2][18] , \ADDER_IN_from_sum[2][17] , 
        \ADDER_IN_from_sum[2][16] , \ADDER_IN_from_sum[2][15] , 
        \ADDER_IN_from_sum[2][14] , \ADDER_IN_from_sum[2][13] , 
        \ADDER_IN_from_sum[2][12] , \ADDER_IN_from_sum[2][11] , 
        \ADDER_IN_from_sum[2][10] , \ADDER_IN_from_sum[2][9] , 
        \ADDER_IN_from_sum[2][8] , \ADDER_IN_from_sum[2][7] , 
        \ADDER_IN_from_sum[2][6] , \ADDER_IN_from_sum[2][5] , 
        \ADDER_IN_from_sum[2][4] , \ADDER_IN_from_sum[2][3] , 
        \ADDER_IN_from_sum[2][2] , \ADDER_IN_from_sum[2][1] , 
        \ADDER_IN_from_sum[2][0] }), .B({\ADDER_IN_from_mux[4][63] , 
        \ADDER_IN_from_mux[4][62] , \ADDER_IN_from_mux[4][61] , 
        \ADDER_IN_from_mux[4][60] , \ADDER_IN_from_mux[4][59] , 
        \ADDER_IN_from_mux[4][58] , \ADDER_IN_from_mux[4][57] , 
        \ADDER_IN_from_mux[4][56] , \ADDER_IN_from_mux[4][55] , 
        \ADDER_IN_from_mux[4][54] , \ADDER_IN_from_mux[4][53] , 
        \ADDER_IN_from_mux[4][52] , \ADDER_IN_from_mux[4][51] , 
        \ADDER_IN_from_mux[4][50] , \ADDER_IN_from_mux[4][49] , 
        \ADDER_IN_from_mux[4][48] , \ADDER_IN_from_mux[4][47] , 
        \ADDER_IN_from_mux[4][46] , \ADDER_IN_from_mux[4][45] , 
        \ADDER_IN_from_mux[4][44] , \ADDER_IN_from_mux[4][43] , 
        \ADDER_IN_from_mux[4][42] , \ADDER_IN_from_mux[4][41] , 
        \ADDER_IN_from_mux[4][40] , \ADDER_IN_from_mux[4][39] , 
        \ADDER_IN_from_mux[4][38] , \ADDER_IN_from_mux[4][37] , 
        \ADDER_IN_from_mux[4][36] , \ADDER_IN_from_mux[4][35] , 
        \ADDER_IN_from_mux[4][34] , \ADDER_IN_from_mux[4][33] , 
        \ADDER_IN_from_mux[4][32] , \ADDER_IN_from_mux[4][31] , 
        \ADDER_IN_from_mux[4][30] , \ADDER_IN_from_mux[4][29] , 
        \ADDER_IN_from_mux[4][28] , \ADDER_IN_from_mux[4][27] , 
        \ADDER_IN_from_mux[4][26] , \ADDER_IN_from_mux[4][25] , 
        \ADDER_IN_from_mux[4][24] , \ADDER_IN_from_mux[4][23] , 
        \ADDER_IN_from_mux[4][22] , \ADDER_IN_from_mux[4][21] , 
        \ADDER_IN_from_mux[4][20] , \ADDER_IN_from_mux[4][19] , 
        \ADDER_IN_from_mux[4][18] , \ADDER_IN_from_mux[4][17] , 
        \ADDER_IN_from_mux[4][16] , \ADDER_IN_from_mux[4][15] , 
        \ADDER_IN_from_mux[4][14] , \ADDER_IN_from_mux[4][13] , 
        \ADDER_IN_from_mux[4][12] , \ADDER_IN_from_mux[4][11] , 
        \ADDER_IN_from_mux[4][10] , \ADDER_IN_from_mux[4][9] , 
        \ADDER_IN_from_mux[4][8] , \ADDER_IN_from_mux[4][7] , 
        \ADDER_IN_from_mux[4][6] , \ADDER_IN_from_mux[4][5] , 
        \ADDER_IN_from_mux[4][4] , \ADDER_IN_from_mux[4][3] , 
        \ADDER_IN_from_mux[4][2] , \ADDER_IN_from_mux[4][1] , 
        \ADDER_IN_from_mux[4][0] }), .S({\ADDER_IN_from_sum[3][63] , 
        \ADDER_IN_from_sum[3][62] , \ADDER_IN_from_sum[3][61] , 
        \ADDER_IN_from_sum[3][60] , \ADDER_IN_from_sum[3][59] , 
        \ADDER_IN_from_sum[3][58] , \ADDER_IN_from_sum[3][57] , 
        \ADDER_IN_from_sum[3][56] , \ADDER_IN_from_sum[3][55] , 
        \ADDER_IN_from_sum[3][54] , \ADDER_IN_from_sum[3][53] , 
        \ADDER_IN_from_sum[3][52] , \ADDER_IN_from_sum[3][51] , 
        \ADDER_IN_from_sum[3][50] , \ADDER_IN_from_sum[3][49] , 
        \ADDER_IN_from_sum[3][48] , \ADDER_IN_from_sum[3][47] , 
        \ADDER_IN_from_sum[3][46] , \ADDER_IN_from_sum[3][45] , 
        \ADDER_IN_from_sum[3][44] , \ADDER_IN_from_sum[3][43] , 
        \ADDER_IN_from_sum[3][42] , \ADDER_IN_from_sum[3][41] , 
        \ADDER_IN_from_sum[3][40] , \ADDER_IN_from_sum[3][39] , 
        \ADDER_IN_from_sum[3][38] , \ADDER_IN_from_sum[3][37] , 
        \ADDER_IN_from_sum[3][36] , \ADDER_IN_from_sum[3][35] , 
        \ADDER_IN_from_sum[3][34] , \ADDER_IN_from_sum[3][33] , 
        \ADDER_IN_from_sum[3][32] , \ADDER_IN_from_sum[3][31] , 
        \ADDER_IN_from_sum[3][30] , \ADDER_IN_from_sum[3][29] , 
        \ADDER_IN_from_sum[3][28] , \ADDER_IN_from_sum[3][27] , 
        \ADDER_IN_from_sum[3][26] , \ADDER_IN_from_sum[3][25] , 
        \ADDER_IN_from_sum[3][24] , \ADDER_IN_from_sum[3][23] , 
        \ADDER_IN_from_sum[3][22] , \ADDER_IN_from_sum[3][21] , 
        \ADDER_IN_from_sum[3][20] , \ADDER_IN_from_sum[3][19] , 
        \ADDER_IN_from_sum[3][18] , \ADDER_IN_from_sum[3][17] , 
        \ADDER_IN_from_sum[3][16] , \ADDER_IN_from_sum[3][15] , 
        \ADDER_IN_from_sum[3][14] , \ADDER_IN_from_sum[3][13] , 
        \ADDER_IN_from_sum[3][12] , \ADDER_IN_from_sum[3][11] , 
        \ADDER_IN_from_sum[3][10] , \ADDER_IN_from_sum[3][9] , 
        \ADDER_IN_from_sum[3][8] , \ADDER_IN_from_sum[3][7] , 
        \ADDER_IN_from_sum[3][6] , \ADDER_IN_from_sum[3][5] , 
        \ADDER_IN_from_sum[3][4] , \ADDER_IN_from_sum[3][3] , 
        \ADDER_IN_from_sum[3][2] , \ADDER_IN_from_sum[3][1] , 
        \ADDER_IN_from_sum[3][0] }) );
  RCA_NBIT64_11 RCA_n_3 ( .A({\ADDER_IN_from_sum[3][63] , 
        \ADDER_IN_from_sum[3][62] , \ADDER_IN_from_sum[3][61] , 
        \ADDER_IN_from_sum[3][60] , \ADDER_IN_from_sum[3][59] , 
        \ADDER_IN_from_sum[3][58] , \ADDER_IN_from_sum[3][57] , 
        \ADDER_IN_from_sum[3][56] , \ADDER_IN_from_sum[3][55] , 
        \ADDER_IN_from_sum[3][54] , \ADDER_IN_from_sum[3][53] , 
        \ADDER_IN_from_sum[3][52] , \ADDER_IN_from_sum[3][51] , 
        \ADDER_IN_from_sum[3][50] , \ADDER_IN_from_sum[3][49] , 
        \ADDER_IN_from_sum[3][48] , \ADDER_IN_from_sum[3][47] , 
        \ADDER_IN_from_sum[3][46] , \ADDER_IN_from_sum[3][45] , 
        \ADDER_IN_from_sum[3][44] , \ADDER_IN_from_sum[3][43] , 
        \ADDER_IN_from_sum[3][42] , \ADDER_IN_from_sum[3][41] , 
        \ADDER_IN_from_sum[3][40] , \ADDER_IN_from_sum[3][39] , 
        \ADDER_IN_from_sum[3][38] , \ADDER_IN_from_sum[3][37] , 
        \ADDER_IN_from_sum[3][36] , \ADDER_IN_from_sum[3][35] , 
        \ADDER_IN_from_sum[3][34] , \ADDER_IN_from_sum[3][33] , 
        \ADDER_IN_from_sum[3][32] , \ADDER_IN_from_sum[3][31] , 
        \ADDER_IN_from_sum[3][30] , \ADDER_IN_from_sum[3][29] , 
        \ADDER_IN_from_sum[3][28] , \ADDER_IN_from_sum[3][27] , 
        \ADDER_IN_from_sum[3][26] , \ADDER_IN_from_sum[3][25] , 
        \ADDER_IN_from_sum[3][24] , \ADDER_IN_from_sum[3][23] , 
        \ADDER_IN_from_sum[3][22] , \ADDER_IN_from_sum[3][21] , 
        \ADDER_IN_from_sum[3][20] , \ADDER_IN_from_sum[3][19] , 
        \ADDER_IN_from_sum[3][18] , \ADDER_IN_from_sum[3][17] , 
        \ADDER_IN_from_sum[3][16] , \ADDER_IN_from_sum[3][15] , 
        \ADDER_IN_from_sum[3][14] , \ADDER_IN_from_sum[3][13] , 
        \ADDER_IN_from_sum[3][12] , \ADDER_IN_from_sum[3][11] , 
        \ADDER_IN_from_sum[3][10] , \ADDER_IN_from_sum[3][9] , 
        \ADDER_IN_from_sum[3][8] , \ADDER_IN_from_sum[3][7] , 
        \ADDER_IN_from_sum[3][6] , \ADDER_IN_from_sum[3][5] , 
        \ADDER_IN_from_sum[3][4] , \ADDER_IN_from_sum[3][3] , 
        \ADDER_IN_from_sum[3][2] , \ADDER_IN_from_sum[3][1] , 
        \ADDER_IN_from_sum[3][0] }), .B({\ADDER_IN_from_mux[5][63] , 
        \ADDER_IN_from_mux[5][62] , \ADDER_IN_from_mux[5][61] , 
        \ADDER_IN_from_mux[5][60] , \ADDER_IN_from_mux[5][59] , 
        \ADDER_IN_from_mux[5][58] , \ADDER_IN_from_mux[5][57] , 
        \ADDER_IN_from_mux[5][56] , \ADDER_IN_from_mux[5][55] , 
        \ADDER_IN_from_mux[5][54] , \ADDER_IN_from_mux[5][53] , 
        \ADDER_IN_from_mux[5][52] , \ADDER_IN_from_mux[5][51] , 
        \ADDER_IN_from_mux[5][50] , \ADDER_IN_from_mux[5][49] , 
        \ADDER_IN_from_mux[5][48] , \ADDER_IN_from_mux[5][47] , 
        \ADDER_IN_from_mux[5][46] , \ADDER_IN_from_mux[5][45] , 
        \ADDER_IN_from_mux[5][44] , \ADDER_IN_from_mux[5][43] , 
        \ADDER_IN_from_mux[5][42] , \ADDER_IN_from_mux[5][41] , 
        \ADDER_IN_from_mux[5][40] , \ADDER_IN_from_mux[5][39] , 
        \ADDER_IN_from_mux[5][38] , \ADDER_IN_from_mux[5][37] , 
        \ADDER_IN_from_mux[5][36] , \ADDER_IN_from_mux[5][35] , 
        \ADDER_IN_from_mux[5][34] , \ADDER_IN_from_mux[5][33] , 
        \ADDER_IN_from_mux[5][32] , \ADDER_IN_from_mux[5][31] , 
        \ADDER_IN_from_mux[5][30] , \ADDER_IN_from_mux[5][29] , 
        \ADDER_IN_from_mux[5][28] , \ADDER_IN_from_mux[5][27] , 
        \ADDER_IN_from_mux[5][26] , \ADDER_IN_from_mux[5][25] , 
        \ADDER_IN_from_mux[5][24] , \ADDER_IN_from_mux[5][23] , 
        \ADDER_IN_from_mux[5][22] , \ADDER_IN_from_mux[5][21] , 
        \ADDER_IN_from_mux[5][20] , \ADDER_IN_from_mux[5][19] , 
        \ADDER_IN_from_mux[5][18] , \ADDER_IN_from_mux[5][17] , 
        \ADDER_IN_from_mux[5][16] , \ADDER_IN_from_mux[5][15] , 
        \ADDER_IN_from_mux[5][14] , \ADDER_IN_from_mux[5][13] , 
        \ADDER_IN_from_mux[5][12] , \ADDER_IN_from_mux[5][11] , 
        \ADDER_IN_from_mux[5][10] , \ADDER_IN_from_mux[5][9] , 
        \ADDER_IN_from_mux[5][8] , \ADDER_IN_from_mux[5][7] , 
        \ADDER_IN_from_mux[5][6] , \ADDER_IN_from_mux[5][5] , 
        \ADDER_IN_from_mux[5][4] , \ADDER_IN_from_mux[5][3] , 
        \ADDER_IN_from_mux[5][2] , \ADDER_IN_from_mux[5][1] , 
        \ADDER_IN_from_mux[5][0] }), .S({\ADDER_IN_from_sum[4][63] , 
        \ADDER_IN_from_sum[4][62] , \ADDER_IN_from_sum[4][61] , 
        \ADDER_IN_from_sum[4][60] , \ADDER_IN_from_sum[4][59] , 
        \ADDER_IN_from_sum[4][58] , \ADDER_IN_from_sum[4][57] , 
        \ADDER_IN_from_sum[4][56] , \ADDER_IN_from_sum[4][55] , 
        \ADDER_IN_from_sum[4][54] , \ADDER_IN_from_sum[4][53] , 
        \ADDER_IN_from_sum[4][52] , \ADDER_IN_from_sum[4][51] , 
        \ADDER_IN_from_sum[4][50] , \ADDER_IN_from_sum[4][49] , 
        \ADDER_IN_from_sum[4][48] , \ADDER_IN_from_sum[4][47] , 
        \ADDER_IN_from_sum[4][46] , \ADDER_IN_from_sum[4][45] , 
        \ADDER_IN_from_sum[4][44] , \ADDER_IN_from_sum[4][43] , 
        \ADDER_IN_from_sum[4][42] , \ADDER_IN_from_sum[4][41] , 
        \ADDER_IN_from_sum[4][40] , \ADDER_IN_from_sum[4][39] , 
        \ADDER_IN_from_sum[4][38] , \ADDER_IN_from_sum[4][37] , 
        \ADDER_IN_from_sum[4][36] , \ADDER_IN_from_sum[4][35] , 
        \ADDER_IN_from_sum[4][34] , \ADDER_IN_from_sum[4][33] , 
        \ADDER_IN_from_sum[4][32] , \ADDER_IN_from_sum[4][31] , 
        \ADDER_IN_from_sum[4][30] , \ADDER_IN_from_sum[4][29] , 
        \ADDER_IN_from_sum[4][28] , \ADDER_IN_from_sum[4][27] , 
        \ADDER_IN_from_sum[4][26] , \ADDER_IN_from_sum[4][25] , 
        \ADDER_IN_from_sum[4][24] , \ADDER_IN_from_sum[4][23] , 
        \ADDER_IN_from_sum[4][22] , \ADDER_IN_from_sum[4][21] , 
        \ADDER_IN_from_sum[4][20] , \ADDER_IN_from_sum[4][19] , 
        \ADDER_IN_from_sum[4][18] , \ADDER_IN_from_sum[4][17] , 
        \ADDER_IN_from_sum[4][16] , \ADDER_IN_from_sum[4][15] , 
        \ADDER_IN_from_sum[4][14] , \ADDER_IN_from_sum[4][13] , 
        \ADDER_IN_from_sum[4][12] , \ADDER_IN_from_sum[4][11] , 
        \ADDER_IN_from_sum[4][10] , \ADDER_IN_from_sum[4][9] , 
        \ADDER_IN_from_sum[4][8] , \ADDER_IN_from_sum[4][7] , 
        \ADDER_IN_from_sum[4][6] , \ADDER_IN_from_sum[4][5] , 
        \ADDER_IN_from_sum[4][4] , \ADDER_IN_from_sum[4][3] , 
        \ADDER_IN_from_sum[4][2] , \ADDER_IN_from_sum[4][1] , 
        \ADDER_IN_from_sum[4][0] }) );
  RCA_NBIT64_10 RCA_n_4 ( .A({\ADDER_IN_from_sum[4][63] , 
        \ADDER_IN_from_sum[4][62] , \ADDER_IN_from_sum[4][61] , 
        \ADDER_IN_from_sum[4][60] , \ADDER_IN_from_sum[4][59] , 
        \ADDER_IN_from_sum[4][58] , \ADDER_IN_from_sum[4][57] , 
        \ADDER_IN_from_sum[4][56] , \ADDER_IN_from_sum[4][55] , 
        \ADDER_IN_from_sum[4][54] , \ADDER_IN_from_sum[4][53] , 
        \ADDER_IN_from_sum[4][52] , \ADDER_IN_from_sum[4][51] , 
        \ADDER_IN_from_sum[4][50] , \ADDER_IN_from_sum[4][49] , 
        \ADDER_IN_from_sum[4][48] , \ADDER_IN_from_sum[4][47] , 
        \ADDER_IN_from_sum[4][46] , \ADDER_IN_from_sum[4][45] , 
        \ADDER_IN_from_sum[4][44] , \ADDER_IN_from_sum[4][43] , 
        \ADDER_IN_from_sum[4][42] , \ADDER_IN_from_sum[4][41] , 
        \ADDER_IN_from_sum[4][40] , \ADDER_IN_from_sum[4][39] , 
        \ADDER_IN_from_sum[4][38] , \ADDER_IN_from_sum[4][37] , 
        \ADDER_IN_from_sum[4][36] , \ADDER_IN_from_sum[4][35] , 
        \ADDER_IN_from_sum[4][34] , \ADDER_IN_from_sum[4][33] , 
        \ADDER_IN_from_sum[4][32] , \ADDER_IN_from_sum[4][31] , 
        \ADDER_IN_from_sum[4][30] , \ADDER_IN_from_sum[4][29] , 
        \ADDER_IN_from_sum[4][28] , \ADDER_IN_from_sum[4][27] , 
        \ADDER_IN_from_sum[4][26] , \ADDER_IN_from_sum[4][25] , 
        \ADDER_IN_from_sum[4][24] , \ADDER_IN_from_sum[4][23] , 
        \ADDER_IN_from_sum[4][22] , \ADDER_IN_from_sum[4][21] , 
        \ADDER_IN_from_sum[4][20] , \ADDER_IN_from_sum[4][19] , 
        \ADDER_IN_from_sum[4][18] , \ADDER_IN_from_sum[4][17] , 
        \ADDER_IN_from_sum[4][16] , \ADDER_IN_from_sum[4][15] , 
        \ADDER_IN_from_sum[4][14] , \ADDER_IN_from_sum[4][13] , 
        \ADDER_IN_from_sum[4][12] , \ADDER_IN_from_sum[4][11] , 
        \ADDER_IN_from_sum[4][10] , \ADDER_IN_from_sum[4][9] , 
        \ADDER_IN_from_sum[4][8] , \ADDER_IN_from_sum[4][7] , 
        \ADDER_IN_from_sum[4][6] , \ADDER_IN_from_sum[4][5] , 
        \ADDER_IN_from_sum[4][4] , \ADDER_IN_from_sum[4][3] , 
        \ADDER_IN_from_sum[4][2] , \ADDER_IN_from_sum[4][1] , 
        \ADDER_IN_from_sum[4][0] }), .B({\ADDER_IN_from_mux[6][63] , 
        \ADDER_IN_from_mux[6][62] , \ADDER_IN_from_mux[6][61] , 
        \ADDER_IN_from_mux[6][60] , \ADDER_IN_from_mux[6][59] , 
        \ADDER_IN_from_mux[6][58] , \ADDER_IN_from_mux[6][57] , 
        \ADDER_IN_from_mux[6][56] , \ADDER_IN_from_mux[6][55] , 
        \ADDER_IN_from_mux[6][54] , \ADDER_IN_from_mux[6][53] , 
        \ADDER_IN_from_mux[6][52] , \ADDER_IN_from_mux[6][51] , 
        \ADDER_IN_from_mux[6][50] , \ADDER_IN_from_mux[6][49] , 
        \ADDER_IN_from_mux[6][48] , \ADDER_IN_from_mux[6][47] , 
        \ADDER_IN_from_mux[6][46] , \ADDER_IN_from_mux[6][45] , 
        \ADDER_IN_from_mux[6][44] , \ADDER_IN_from_mux[6][43] , 
        \ADDER_IN_from_mux[6][42] , \ADDER_IN_from_mux[6][41] , 
        \ADDER_IN_from_mux[6][40] , \ADDER_IN_from_mux[6][39] , 
        \ADDER_IN_from_mux[6][38] , \ADDER_IN_from_mux[6][37] , 
        \ADDER_IN_from_mux[6][36] , \ADDER_IN_from_mux[6][35] , 
        \ADDER_IN_from_mux[6][34] , \ADDER_IN_from_mux[6][33] , 
        \ADDER_IN_from_mux[6][32] , \ADDER_IN_from_mux[6][31] , 
        \ADDER_IN_from_mux[6][30] , \ADDER_IN_from_mux[6][29] , 
        \ADDER_IN_from_mux[6][28] , \ADDER_IN_from_mux[6][27] , 
        \ADDER_IN_from_mux[6][26] , \ADDER_IN_from_mux[6][25] , 
        \ADDER_IN_from_mux[6][24] , \ADDER_IN_from_mux[6][23] , 
        \ADDER_IN_from_mux[6][22] , \ADDER_IN_from_mux[6][21] , 
        \ADDER_IN_from_mux[6][20] , \ADDER_IN_from_mux[6][19] , 
        \ADDER_IN_from_mux[6][18] , \ADDER_IN_from_mux[6][17] , 
        \ADDER_IN_from_mux[6][16] , \ADDER_IN_from_mux[6][15] , 
        \ADDER_IN_from_mux[6][14] , \ADDER_IN_from_mux[6][13] , 
        \ADDER_IN_from_mux[6][12] , \ADDER_IN_from_mux[6][11] , 
        \ADDER_IN_from_mux[6][10] , \ADDER_IN_from_mux[6][9] , 
        \ADDER_IN_from_mux[6][8] , \ADDER_IN_from_mux[6][7] , 
        \ADDER_IN_from_mux[6][6] , \ADDER_IN_from_mux[6][5] , 
        \ADDER_IN_from_mux[6][4] , \ADDER_IN_from_mux[6][3] , 
        \ADDER_IN_from_mux[6][2] , \ADDER_IN_from_mux[6][1] , 
        \ADDER_IN_from_mux[6][0] }), .S({\ADDER_IN_from_sum[5][63] , 
        \ADDER_IN_from_sum[5][62] , \ADDER_IN_from_sum[5][61] , 
        \ADDER_IN_from_sum[5][60] , \ADDER_IN_from_sum[5][59] , 
        \ADDER_IN_from_sum[5][58] , \ADDER_IN_from_sum[5][57] , 
        \ADDER_IN_from_sum[5][56] , \ADDER_IN_from_sum[5][55] , 
        \ADDER_IN_from_sum[5][54] , \ADDER_IN_from_sum[5][53] , 
        \ADDER_IN_from_sum[5][52] , \ADDER_IN_from_sum[5][51] , 
        \ADDER_IN_from_sum[5][50] , \ADDER_IN_from_sum[5][49] , 
        \ADDER_IN_from_sum[5][48] , \ADDER_IN_from_sum[5][47] , 
        \ADDER_IN_from_sum[5][46] , \ADDER_IN_from_sum[5][45] , 
        \ADDER_IN_from_sum[5][44] , \ADDER_IN_from_sum[5][43] , 
        \ADDER_IN_from_sum[5][42] , \ADDER_IN_from_sum[5][41] , 
        \ADDER_IN_from_sum[5][40] , \ADDER_IN_from_sum[5][39] , 
        \ADDER_IN_from_sum[5][38] , \ADDER_IN_from_sum[5][37] , 
        \ADDER_IN_from_sum[5][36] , \ADDER_IN_from_sum[5][35] , 
        \ADDER_IN_from_sum[5][34] , \ADDER_IN_from_sum[5][33] , 
        \ADDER_IN_from_sum[5][32] , \ADDER_IN_from_sum[5][31] , 
        \ADDER_IN_from_sum[5][30] , \ADDER_IN_from_sum[5][29] , 
        \ADDER_IN_from_sum[5][28] , \ADDER_IN_from_sum[5][27] , 
        \ADDER_IN_from_sum[5][26] , \ADDER_IN_from_sum[5][25] , 
        \ADDER_IN_from_sum[5][24] , \ADDER_IN_from_sum[5][23] , 
        \ADDER_IN_from_sum[5][22] , \ADDER_IN_from_sum[5][21] , 
        \ADDER_IN_from_sum[5][20] , \ADDER_IN_from_sum[5][19] , 
        \ADDER_IN_from_sum[5][18] , \ADDER_IN_from_sum[5][17] , 
        \ADDER_IN_from_sum[5][16] , \ADDER_IN_from_sum[5][15] , 
        \ADDER_IN_from_sum[5][14] , \ADDER_IN_from_sum[5][13] , 
        \ADDER_IN_from_sum[5][12] , \ADDER_IN_from_sum[5][11] , 
        \ADDER_IN_from_sum[5][10] , \ADDER_IN_from_sum[5][9] , 
        \ADDER_IN_from_sum[5][8] , \ADDER_IN_from_sum[5][7] , 
        \ADDER_IN_from_sum[5][6] , \ADDER_IN_from_sum[5][5] , 
        \ADDER_IN_from_sum[5][4] , \ADDER_IN_from_sum[5][3] , 
        \ADDER_IN_from_sum[5][2] , \ADDER_IN_from_sum[5][1] , 
        \ADDER_IN_from_sum[5][0] }) );
  RCA_NBIT64_9 RCA_n_5 ( .A({\ADDER_IN_from_sum[5][63] , 
        \ADDER_IN_from_sum[5][62] , \ADDER_IN_from_sum[5][61] , 
        \ADDER_IN_from_sum[5][60] , \ADDER_IN_from_sum[5][59] , 
        \ADDER_IN_from_sum[5][58] , \ADDER_IN_from_sum[5][57] , 
        \ADDER_IN_from_sum[5][56] , \ADDER_IN_from_sum[5][55] , 
        \ADDER_IN_from_sum[5][54] , \ADDER_IN_from_sum[5][53] , 
        \ADDER_IN_from_sum[5][52] , \ADDER_IN_from_sum[5][51] , 
        \ADDER_IN_from_sum[5][50] , \ADDER_IN_from_sum[5][49] , 
        \ADDER_IN_from_sum[5][48] , \ADDER_IN_from_sum[5][47] , 
        \ADDER_IN_from_sum[5][46] , \ADDER_IN_from_sum[5][45] , 
        \ADDER_IN_from_sum[5][44] , \ADDER_IN_from_sum[5][43] , 
        \ADDER_IN_from_sum[5][42] , \ADDER_IN_from_sum[5][41] , 
        \ADDER_IN_from_sum[5][40] , \ADDER_IN_from_sum[5][39] , 
        \ADDER_IN_from_sum[5][38] , \ADDER_IN_from_sum[5][37] , 
        \ADDER_IN_from_sum[5][36] , \ADDER_IN_from_sum[5][35] , 
        \ADDER_IN_from_sum[5][34] , \ADDER_IN_from_sum[5][33] , 
        \ADDER_IN_from_sum[5][32] , \ADDER_IN_from_sum[5][31] , 
        \ADDER_IN_from_sum[5][30] , \ADDER_IN_from_sum[5][29] , 
        \ADDER_IN_from_sum[5][28] , \ADDER_IN_from_sum[5][27] , 
        \ADDER_IN_from_sum[5][26] , \ADDER_IN_from_sum[5][25] , 
        \ADDER_IN_from_sum[5][24] , \ADDER_IN_from_sum[5][23] , 
        \ADDER_IN_from_sum[5][22] , \ADDER_IN_from_sum[5][21] , 
        \ADDER_IN_from_sum[5][20] , \ADDER_IN_from_sum[5][19] , 
        \ADDER_IN_from_sum[5][18] , \ADDER_IN_from_sum[5][17] , 
        \ADDER_IN_from_sum[5][16] , \ADDER_IN_from_sum[5][15] , 
        \ADDER_IN_from_sum[5][14] , \ADDER_IN_from_sum[5][13] , 
        \ADDER_IN_from_sum[5][12] , \ADDER_IN_from_sum[5][11] , 
        \ADDER_IN_from_sum[5][10] , \ADDER_IN_from_sum[5][9] , 
        \ADDER_IN_from_sum[5][8] , \ADDER_IN_from_sum[5][7] , 
        \ADDER_IN_from_sum[5][6] , \ADDER_IN_from_sum[5][5] , 
        \ADDER_IN_from_sum[5][4] , \ADDER_IN_from_sum[5][3] , 
        \ADDER_IN_from_sum[5][2] , \ADDER_IN_from_sum[5][1] , 
        \ADDER_IN_from_sum[5][0] }), .B({\ADDER_IN_from_mux[7][63] , 
        \ADDER_IN_from_mux[7][62] , \ADDER_IN_from_mux[7][61] , 
        \ADDER_IN_from_mux[7][60] , \ADDER_IN_from_mux[7][59] , 
        \ADDER_IN_from_mux[7][58] , \ADDER_IN_from_mux[7][57] , 
        \ADDER_IN_from_mux[7][56] , \ADDER_IN_from_mux[7][55] , 
        \ADDER_IN_from_mux[7][54] , \ADDER_IN_from_mux[7][53] , 
        \ADDER_IN_from_mux[7][52] , \ADDER_IN_from_mux[7][51] , 
        \ADDER_IN_from_mux[7][50] , \ADDER_IN_from_mux[7][49] , 
        \ADDER_IN_from_mux[7][48] , \ADDER_IN_from_mux[7][47] , 
        \ADDER_IN_from_mux[7][46] , \ADDER_IN_from_mux[7][45] , 
        \ADDER_IN_from_mux[7][44] , \ADDER_IN_from_mux[7][43] , 
        \ADDER_IN_from_mux[7][42] , \ADDER_IN_from_mux[7][41] , 
        \ADDER_IN_from_mux[7][40] , \ADDER_IN_from_mux[7][39] , 
        \ADDER_IN_from_mux[7][38] , \ADDER_IN_from_mux[7][37] , 
        \ADDER_IN_from_mux[7][36] , \ADDER_IN_from_mux[7][35] , 
        \ADDER_IN_from_mux[7][34] , \ADDER_IN_from_mux[7][33] , 
        \ADDER_IN_from_mux[7][32] , \ADDER_IN_from_mux[7][31] , 
        \ADDER_IN_from_mux[7][30] , \ADDER_IN_from_mux[7][29] , 
        \ADDER_IN_from_mux[7][28] , \ADDER_IN_from_mux[7][27] , 
        \ADDER_IN_from_mux[7][26] , \ADDER_IN_from_mux[7][25] , 
        \ADDER_IN_from_mux[7][24] , \ADDER_IN_from_mux[7][23] , 
        \ADDER_IN_from_mux[7][22] , \ADDER_IN_from_mux[7][21] , 
        \ADDER_IN_from_mux[7][20] , \ADDER_IN_from_mux[7][19] , 
        \ADDER_IN_from_mux[7][18] , \ADDER_IN_from_mux[7][17] , 
        \ADDER_IN_from_mux[7][16] , \ADDER_IN_from_mux[7][15] , 
        \ADDER_IN_from_mux[7][14] , \ADDER_IN_from_mux[7][13] , 
        \ADDER_IN_from_mux[7][12] , \ADDER_IN_from_mux[7][11] , 
        \ADDER_IN_from_mux[7][10] , \ADDER_IN_from_mux[7][9] , 
        \ADDER_IN_from_mux[7][8] , \ADDER_IN_from_mux[7][7] , 
        \ADDER_IN_from_mux[7][6] , \ADDER_IN_from_mux[7][5] , 
        \ADDER_IN_from_mux[7][4] , \ADDER_IN_from_mux[7][3] , 
        \ADDER_IN_from_mux[7][2] , \ADDER_IN_from_mux[7][1] , 
        \ADDER_IN_from_mux[7][0] }), .S({\ADDER_IN_from_sum[6][63] , 
        \ADDER_IN_from_sum[6][62] , \ADDER_IN_from_sum[6][61] , 
        \ADDER_IN_from_sum[6][60] , \ADDER_IN_from_sum[6][59] , 
        \ADDER_IN_from_sum[6][58] , \ADDER_IN_from_sum[6][57] , 
        \ADDER_IN_from_sum[6][56] , \ADDER_IN_from_sum[6][55] , 
        \ADDER_IN_from_sum[6][54] , \ADDER_IN_from_sum[6][53] , 
        \ADDER_IN_from_sum[6][52] , \ADDER_IN_from_sum[6][51] , 
        \ADDER_IN_from_sum[6][50] , \ADDER_IN_from_sum[6][49] , 
        \ADDER_IN_from_sum[6][48] , \ADDER_IN_from_sum[6][47] , 
        \ADDER_IN_from_sum[6][46] , \ADDER_IN_from_sum[6][45] , 
        \ADDER_IN_from_sum[6][44] , \ADDER_IN_from_sum[6][43] , 
        \ADDER_IN_from_sum[6][42] , \ADDER_IN_from_sum[6][41] , 
        \ADDER_IN_from_sum[6][40] , \ADDER_IN_from_sum[6][39] , 
        \ADDER_IN_from_sum[6][38] , \ADDER_IN_from_sum[6][37] , 
        \ADDER_IN_from_sum[6][36] , \ADDER_IN_from_sum[6][35] , 
        \ADDER_IN_from_sum[6][34] , \ADDER_IN_from_sum[6][33] , 
        \ADDER_IN_from_sum[6][32] , \ADDER_IN_from_sum[6][31] , 
        \ADDER_IN_from_sum[6][30] , \ADDER_IN_from_sum[6][29] , 
        \ADDER_IN_from_sum[6][28] , \ADDER_IN_from_sum[6][27] , 
        \ADDER_IN_from_sum[6][26] , \ADDER_IN_from_sum[6][25] , 
        \ADDER_IN_from_sum[6][24] , \ADDER_IN_from_sum[6][23] , 
        \ADDER_IN_from_sum[6][22] , \ADDER_IN_from_sum[6][21] , 
        \ADDER_IN_from_sum[6][20] , \ADDER_IN_from_sum[6][19] , 
        \ADDER_IN_from_sum[6][18] , \ADDER_IN_from_sum[6][17] , 
        \ADDER_IN_from_sum[6][16] , \ADDER_IN_from_sum[6][15] , 
        \ADDER_IN_from_sum[6][14] , \ADDER_IN_from_sum[6][13] , 
        \ADDER_IN_from_sum[6][12] , \ADDER_IN_from_sum[6][11] , 
        \ADDER_IN_from_sum[6][10] , \ADDER_IN_from_sum[6][9] , 
        \ADDER_IN_from_sum[6][8] , \ADDER_IN_from_sum[6][7] , 
        \ADDER_IN_from_sum[6][6] , \ADDER_IN_from_sum[6][5] , 
        \ADDER_IN_from_sum[6][4] , \ADDER_IN_from_sum[6][3] , 
        \ADDER_IN_from_sum[6][2] , \ADDER_IN_from_sum[6][1] , 
        \ADDER_IN_from_sum[6][0] }) );
  RCA_NBIT64_8 RCA_n_6 ( .A({\ADDER_IN_from_sum[6][63] , 
        \ADDER_IN_from_sum[6][62] , \ADDER_IN_from_sum[6][61] , 
        \ADDER_IN_from_sum[6][60] , \ADDER_IN_from_sum[6][59] , 
        \ADDER_IN_from_sum[6][58] , \ADDER_IN_from_sum[6][57] , 
        \ADDER_IN_from_sum[6][56] , \ADDER_IN_from_sum[6][55] , 
        \ADDER_IN_from_sum[6][54] , \ADDER_IN_from_sum[6][53] , 
        \ADDER_IN_from_sum[6][52] , \ADDER_IN_from_sum[6][51] , 
        \ADDER_IN_from_sum[6][50] , \ADDER_IN_from_sum[6][49] , 
        \ADDER_IN_from_sum[6][48] , \ADDER_IN_from_sum[6][47] , 
        \ADDER_IN_from_sum[6][46] , \ADDER_IN_from_sum[6][45] , 
        \ADDER_IN_from_sum[6][44] , \ADDER_IN_from_sum[6][43] , 
        \ADDER_IN_from_sum[6][42] , \ADDER_IN_from_sum[6][41] , 
        \ADDER_IN_from_sum[6][40] , \ADDER_IN_from_sum[6][39] , 
        \ADDER_IN_from_sum[6][38] , \ADDER_IN_from_sum[6][37] , 
        \ADDER_IN_from_sum[6][36] , \ADDER_IN_from_sum[6][35] , 
        \ADDER_IN_from_sum[6][34] , \ADDER_IN_from_sum[6][33] , 
        \ADDER_IN_from_sum[6][32] , \ADDER_IN_from_sum[6][31] , 
        \ADDER_IN_from_sum[6][30] , \ADDER_IN_from_sum[6][29] , 
        \ADDER_IN_from_sum[6][28] , \ADDER_IN_from_sum[6][27] , 
        \ADDER_IN_from_sum[6][26] , \ADDER_IN_from_sum[6][25] , 
        \ADDER_IN_from_sum[6][24] , \ADDER_IN_from_sum[6][23] , 
        \ADDER_IN_from_sum[6][22] , \ADDER_IN_from_sum[6][21] , 
        \ADDER_IN_from_sum[6][20] , \ADDER_IN_from_sum[6][19] , 
        \ADDER_IN_from_sum[6][18] , \ADDER_IN_from_sum[6][17] , 
        \ADDER_IN_from_sum[6][16] , \ADDER_IN_from_sum[6][15] , 
        \ADDER_IN_from_sum[6][14] , \ADDER_IN_from_sum[6][13] , 
        \ADDER_IN_from_sum[6][12] , \ADDER_IN_from_sum[6][11] , 
        \ADDER_IN_from_sum[6][10] , \ADDER_IN_from_sum[6][9] , 
        \ADDER_IN_from_sum[6][8] , \ADDER_IN_from_sum[6][7] , 
        \ADDER_IN_from_sum[6][6] , \ADDER_IN_from_sum[6][5] , 
        \ADDER_IN_from_sum[6][4] , \ADDER_IN_from_sum[6][3] , 
        \ADDER_IN_from_sum[6][2] , \ADDER_IN_from_sum[6][1] , 
        \ADDER_IN_from_sum[6][0] }), .B({\ADDER_IN_from_mux[8][63] , 
        \ADDER_IN_from_mux[8][62] , \ADDER_IN_from_mux[8][61] , 
        \ADDER_IN_from_mux[8][60] , \ADDER_IN_from_mux[8][59] , 
        \ADDER_IN_from_mux[8][58] , \ADDER_IN_from_mux[8][57] , 
        \ADDER_IN_from_mux[8][56] , \ADDER_IN_from_mux[8][55] , 
        \ADDER_IN_from_mux[8][54] , \ADDER_IN_from_mux[8][53] , 
        \ADDER_IN_from_mux[8][52] , \ADDER_IN_from_mux[8][51] , 
        \ADDER_IN_from_mux[8][50] , \ADDER_IN_from_mux[8][49] , 
        \ADDER_IN_from_mux[8][48] , \ADDER_IN_from_mux[8][47] , 
        \ADDER_IN_from_mux[8][46] , \ADDER_IN_from_mux[8][45] , 
        \ADDER_IN_from_mux[8][44] , \ADDER_IN_from_mux[8][43] , 
        \ADDER_IN_from_mux[8][42] , \ADDER_IN_from_mux[8][41] , 
        \ADDER_IN_from_mux[8][40] , \ADDER_IN_from_mux[8][39] , 
        \ADDER_IN_from_mux[8][38] , \ADDER_IN_from_mux[8][37] , 
        \ADDER_IN_from_mux[8][36] , \ADDER_IN_from_mux[8][35] , 
        \ADDER_IN_from_mux[8][34] , \ADDER_IN_from_mux[8][33] , 
        \ADDER_IN_from_mux[8][32] , \ADDER_IN_from_mux[8][31] , 
        \ADDER_IN_from_mux[8][30] , \ADDER_IN_from_mux[8][29] , 
        \ADDER_IN_from_mux[8][28] , \ADDER_IN_from_mux[8][27] , 
        \ADDER_IN_from_mux[8][26] , \ADDER_IN_from_mux[8][25] , 
        \ADDER_IN_from_mux[8][24] , \ADDER_IN_from_mux[8][23] , 
        \ADDER_IN_from_mux[8][22] , \ADDER_IN_from_mux[8][21] , 
        \ADDER_IN_from_mux[8][20] , \ADDER_IN_from_mux[8][19] , 
        \ADDER_IN_from_mux[8][18] , \ADDER_IN_from_mux[8][17] , 
        \ADDER_IN_from_mux[8][16] , \ADDER_IN_from_mux[8][15] , 
        \ADDER_IN_from_mux[8][14] , \ADDER_IN_from_mux[8][13] , 
        \ADDER_IN_from_mux[8][12] , \ADDER_IN_from_mux[8][11] , 
        \ADDER_IN_from_mux[8][10] , \ADDER_IN_from_mux[8][9] , 
        \ADDER_IN_from_mux[8][8] , \ADDER_IN_from_mux[8][7] , 
        \ADDER_IN_from_mux[8][6] , \ADDER_IN_from_mux[8][5] , 
        \ADDER_IN_from_mux[8][4] , \ADDER_IN_from_mux[8][3] , 
        \ADDER_IN_from_mux[8][2] , \ADDER_IN_from_mux[8][1] , 
        \ADDER_IN_from_mux[8][0] }), .S({\ADDER_IN_from_sum[7][63] , 
        \ADDER_IN_from_sum[7][62] , \ADDER_IN_from_sum[7][61] , 
        \ADDER_IN_from_sum[7][60] , \ADDER_IN_from_sum[7][59] , 
        \ADDER_IN_from_sum[7][58] , \ADDER_IN_from_sum[7][57] , 
        \ADDER_IN_from_sum[7][56] , \ADDER_IN_from_sum[7][55] , 
        \ADDER_IN_from_sum[7][54] , \ADDER_IN_from_sum[7][53] , 
        \ADDER_IN_from_sum[7][52] , \ADDER_IN_from_sum[7][51] , 
        \ADDER_IN_from_sum[7][50] , \ADDER_IN_from_sum[7][49] , 
        \ADDER_IN_from_sum[7][48] , \ADDER_IN_from_sum[7][47] , 
        \ADDER_IN_from_sum[7][46] , \ADDER_IN_from_sum[7][45] , 
        \ADDER_IN_from_sum[7][44] , \ADDER_IN_from_sum[7][43] , 
        \ADDER_IN_from_sum[7][42] , \ADDER_IN_from_sum[7][41] , 
        \ADDER_IN_from_sum[7][40] , \ADDER_IN_from_sum[7][39] , 
        \ADDER_IN_from_sum[7][38] , \ADDER_IN_from_sum[7][37] , 
        \ADDER_IN_from_sum[7][36] , \ADDER_IN_from_sum[7][35] , 
        \ADDER_IN_from_sum[7][34] , \ADDER_IN_from_sum[7][33] , 
        \ADDER_IN_from_sum[7][32] , \ADDER_IN_from_sum[7][31] , 
        \ADDER_IN_from_sum[7][30] , \ADDER_IN_from_sum[7][29] , 
        \ADDER_IN_from_sum[7][28] , \ADDER_IN_from_sum[7][27] , 
        \ADDER_IN_from_sum[7][26] , \ADDER_IN_from_sum[7][25] , 
        \ADDER_IN_from_sum[7][24] , \ADDER_IN_from_sum[7][23] , 
        \ADDER_IN_from_sum[7][22] , \ADDER_IN_from_sum[7][21] , 
        \ADDER_IN_from_sum[7][20] , \ADDER_IN_from_sum[7][19] , 
        \ADDER_IN_from_sum[7][18] , \ADDER_IN_from_sum[7][17] , 
        \ADDER_IN_from_sum[7][16] , \ADDER_IN_from_sum[7][15] , 
        \ADDER_IN_from_sum[7][14] , \ADDER_IN_from_sum[7][13] , 
        \ADDER_IN_from_sum[7][12] , \ADDER_IN_from_sum[7][11] , 
        \ADDER_IN_from_sum[7][10] , \ADDER_IN_from_sum[7][9] , 
        \ADDER_IN_from_sum[7][8] , \ADDER_IN_from_sum[7][7] , 
        \ADDER_IN_from_sum[7][6] , \ADDER_IN_from_sum[7][5] , 
        \ADDER_IN_from_sum[7][4] , \ADDER_IN_from_sum[7][3] , 
        \ADDER_IN_from_sum[7][2] , \ADDER_IN_from_sum[7][1] , 
        \ADDER_IN_from_sum[7][0] }) );
  RCA_NBIT64_7 RCA_n_7 ( .A({\ADDER_IN_from_sum[7][63] , 
        \ADDER_IN_from_sum[7][62] , \ADDER_IN_from_sum[7][61] , 
        \ADDER_IN_from_sum[7][60] , \ADDER_IN_from_sum[7][59] , 
        \ADDER_IN_from_sum[7][58] , \ADDER_IN_from_sum[7][57] , 
        \ADDER_IN_from_sum[7][56] , \ADDER_IN_from_sum[7][55] , 
        \ADDER_IN_from_sum[7][54] , \ADDER_IN_from_sum[7][53] , 
        \ADDER_IN_from_sum[7][52] , \ADDER_IN_from_sum[7][51] , 
        \ADDER_IN_from_sum[7][50] , \ADDER_IN_from_sum[7][49] , 
        \ADDER_IN_from_sum[7][48] , \ADDER_IN_from_sum[7][47] , 
        \ADDER_IN_from_sum[7][46] , \ADDER_IN_from_sum[7][45] , 
        \ADDER_IN_from_sum[7][44] , \ADDER_IN_from_sum[7][43] , 
        \ADDER_IN_from_sum[7][42] , \ADDER_IN_from_sum[7][41] , 
        \ADDER_IN_from_sum[7][40] , \ADDER_IN_from_sum[7][39] , 
        \ADDER_IN_from_sum[7][38] , \ADDER_IN_from_sum[7][37] , 
        \ADDER_IN_from_sum[7][36] , \ADDER_IN_from_sum[7][35] , 
        \ADDER_IN_from_sum[7][34] , \ADDER_IN_from_sum[7][33] , 
        \ADDER_IN_from_sum[7][32] , \ADDER_IN_from_sum[7][31] , 
        \ADDER_IN_from_sum[7][30] , \ADDER_IN_from_sum[7][29] , 
        \ADDER_IN_from_sum[7][28] , \ADDER_IN_from_sum[7][27] , 
        \ADDER_IN_from_sum[7][26] , \ADDER_IN_from_sum[7][25] , 
        \ADDER_IN_from_sum[7][24] , \ADDER_IN_from_sum[7][23] , 
        \ADDER_IN_from_sum[7][22] , \ADDER_IN_from_sum[7][21] , 
        \ADDER_IN_from_sum[7][20] , \ADDER_IN_from_sum[7][19] , 
        \ADDER_IN_from_sum[7][18] , \ADDER_IN_from_sum[7][17] , 
        \ADDER_IN_from_sum[7][16] , \ADDER_IN_from_sum[7][15] , 
        \ADDER_IN_from_sum[7][14] , \ADDER_IN_from_sum[7][13] , 
        \ADDER_IN_from_sum[7][12] , \ADDER_IN_from_sum[7][11] , 
        \ADDER_IN_from_sum[7][10] , \ADDER_IN_from_sum[7][9] , 
        \ADDER_IN_from_sum[7][8] , \ADDER_IN_from_sum[7][7] , 
        \ADDER_IN_from_sum[7][6] , \ADDER_IN_from_sum[7][5] , 
        \ADDER_IN_from_sum[7][4] , \ADDER_IN_from_sum[7][3] , 
        \ADDER_IN_from_sum[7][2] , \ADDER_IN_from_sum[7][1] , 
        \ADDER_IN_from_sum[7][0] }), .B({\ADDER_IN_from_mux[9][63] , 
        \ADDER_IN_from_mux[9][62] , \ADDER_IN_from_mux[9][61] , 
        \ADDER_IN_from_mux[9][60] , \ADDER_IN_from_mux[9][59] , 
        \ADDER_IN_from_mux[9][58] , \ADDER_IN_from_mux[9][57] , 
        \ADDER_IN_from_mux[9][56] , \ADDER_IN_from_mux[9][55] , 
        \ADDER_IN_from_mux[9][54] , \ADDER_IN_from_mux[9][53] , 
        \ADDER_IN_from_mux[9][52] , \ADDER_IN_from_mux[9][51] , 
        \ADDER_IN_from_mux[9][50] , \ADDER_IN_from_mux[9][49] , 
        \ADDER_IN_from_mux[9][48] , \ADDER_IN_from_mux[9][47] , 
        \ADDER_IN_from_mux[9][46] , \ADDER_IN_from_mux[9][45] , 
        \ADDER_IN_from_mux[9][44] , \ADDER_IN_from_mux[9][43] , 
        \ADDER_IN_from_mux[9][42] , \ADDER_IN_from_mux[9][41] , 
        \ADDER_IN_from_mux[9][40] , \ADDER_IN_from_mux[9][39] , 
        \ADDER_IN_from_mux[9][38] , \ADDER_IN_from_mux[9][37] , 
        \ADDER_IN_from_mux[9][36] , \ADDER_IN_from_mux[9][35] , 
        \ADDER_IN_from_mux[9][34] , \ADDER_IN_from_mux[9][33] , 
        \ADDER_IN_from_mux[9][32] , \ADDER_IN_from_mux[9][31] , 
        \ADDER_IN_from_mux[9][30] , \ADDER_IN_from_mux[9][29] , 
        \ADDER_IN_from_mux[9][28] , \ADDER_IN_from_mux[9][27] , 
        \ADDER_IN_from_mux[9][26] , \ADDER_IN_from_mux[9][25] , 
        \ADDER_IN_from_mux[9][24] , \ADDER_IN_from_mux[9][23] , 
        \ADDER_IN_from_mux[9][22] , \ADDER_IN_from_mux[9][21] , 
        \ADDER_IN_from_mux[9][20] , \ADDER_IN_from_mux[9][19] , 
        \ADDER_IN_from_mux[9][18] , \ADDER_IN_from_mux[9][17] , 
        \ADDER_IN_from_mux[9][16] , \ADDER_IN_from_mux[9][15] , 
        \ADDER_IN_from_mux[9][14] , \ADDER_IN_from_mux[9][13] , 
        \ADDER_IN_from_mux[9][12] , \ADDER_IN_from_mux[9][11] , 
        \ADDER_IN_from_mux[9][10] , \ADDER_IN_from_mux[9][9] , 
        \ADDER_IN_from_mux[9][8] , \ADDER_IN_from_mux[9][7] , 
        \ADDER_IN_from_mux[9][6] , \ADDER_IN_from_mux[9][5] , 
        \ADDER_IN_from_mux[9][4] , \ADDER_IN_from_mux[9][3] , 
        \ADDER_IN_from_mux[9][2] , \ADDER_IN_from_mux[9][1] , 
        \ADDER_IN_from_mux[9][0] }), .S({\ADDER_IN_from_sum[8][63] , 
        \ADDER_IN_from_sum[8][62] , \ADDER_IN_from_sum[8][61] , 
        \ADDER_IN_from_sum[8][60] , \ADDER_IN_from_sum[8][59] , 
        \ADDER_IN_from_sum[8][58] , \ADDER_IN_from_sum[8][57] , 
        \ADDER_IN_from_sum[8][56] , \ADDER_IN_from_sum[8][55] , 
        \ADDER_IN_from_sum[8][54] , \ADDER_IN_from_sum[8][53] , 
        \ADDER_IN_from_sum[8][52] , \ADDER_IN_from_sum[8][51] , 
        \ADDER_IN_from_sum[8][50] , \ADDER_IN_from_sum[8][49] , 
        \ADDER_IN_from_sum[8][48] , \ADDER_IN_from_sum[8][47] , 
        \ADDER_IN_from_sum[8][46] , \ADDER_IN_from_sum[8][45] , 
        \ADDER_IN_from_sum[8][44] , \ADDER_IN_from_sum[8][43] , 
        \ADDER_IN_from_sum[8][42] , \ADDER_IN_from_sum[8][41] , 
        \ADDER_IN_from_sum[8][40] , \ADDER_IN_from_sum[8][39] , 
        \ADDER_IN_from_sum[8][38] , \ADDER_IN_from_sum[8][37] , 
        \ADDER_IN_from_sum[8][36] , \ADDER_IN_from_sum[8][35] , 
        \ADDER_IN_from_sum[8][34] , \ADDER_IN_from_sum[8][33] , 
        \ADDER_IN_from_sum[8][32] , \ADDER_IN_from_sum[8][31] , 
        \ADDER_IN_from_sum[8][30] , \ADDER_IN_from_sum[8][29] , 
        \ADDER_IN_from_sum[8][28] , \ADDER_IN_from_sum[8][27] , 
        \ADDER_IN_from_sum[8][26] , \ADDER_IN_from_sum[8][25] , 
        \ADDER_IN_from_sum[8][24] , \ADDER_IN_from_sum[8][23] , 
        \ADDER_IN_from_sum[8][22] , \ADDER_IN_from_sum[8][21] , 
        \ADDER_IN_from_sum[8][20] , \ADDER_IN_from_sum[8][19] , 
        \ADDER_IN_from_sum[8][18] , \ADDER_IN_from_sum[8][17] , 
        \ADDER_IN_from_sum[8][16] , \ADDER_IN_from_sum[8][15] , 
        \ADDER_IN_from_sum[8][14] , \ADDER_IN_from_sum[8][13] , 
        \ADDER_IN_from_sum[8][12] , \ADDER_IN_from_sum[8][11] , 
        \ADDER_IN_from_sum[8][10] , \ADDER_IN_from_sum[8][9] , 
        \ADDER_IN_from_sum[8][8] , \ADDER_IN_from_sum[8][7] , 
        \ADDER_IN_from_sum[8][6] , \ADDER_IN_from_sum[8][5] , 
        \ADDER_IN_from_sum[8][4] , \ADDER_IN_from_sum[8][3] , 
        \ADDER_IN_from_sum[8][2] , \ADDER_IN_from_sum[8][1] , 
        \ADDER_IN_from_sum[8][0] }) );
  RCA_NBIT64_6 RCA_n_8 ( .A({\ADDER_IN_from_sum[8][63] , 
        \ADDER_IN_from_sum[8][62] , \ADDER_IN_from_sum[8][61] , 
        \ADDER_IN_from_sum[8][60] , \ADDER_IN_from_sum[8][59] , 
        \ADDER_IN_from_sum[8][58] , \ADDER_IN_from_sum[8][57] , 
        \ADDER_IN_from_sum[8][56] , \ADDER_IN_from_sum[8][55] , 
        \ADDER_IN_from_sum[8][54] , \ADDER_IN_from_sum[8][53] , 
        \ADDER_IN_from_sum[8][52] , \ADDER_IN_from_sum[8][51] , 
        \ADDER_IN_from_sum[8][50] , \ADDER_IN_from_sum[8][49] , 
        \ADDER_IN_from_sum[8][48] , \ADDER_IN_from_sum[8][47] , 
        \ADDER_IN_from_sum[8][46] , \ADDER_IN_from_sum[8][45] , 
        \ADDER_IN_from_sum[8][44] , \ADDER_IN_from_sum[8][43] , 
        \ADDER_IN_from_sum[8][42] , \ADDER_IN_from_sum[8][41] , 
        \ADDER_IN_from_sum[8][40] , \ADDER_IN_from_sum[8][39] , 
        \ADDER_IN_from_sum[8][38] , \ADDER_IN_from_sum[8][37] , 
        \ADDER_IN_from_sum[8][36] , \ADDER_IN_from_sum[8][35] , 
        \ADDER_IN_from_sum[8][34] , \ADDER_IN_from_sum[8][33] , 
        \ADDER_IN_from_sum[8][32] , \ADDER_IN_from_sum[8][31] , 
        \ADDER_IN_from_sum[8][30] , \ADDER_IN_from_sum[8][29] , 
        \ADDER_IN_from_sum[8][28] , \ADDER_IN_from_sum[8][27] , 
        \ADDER_IN_from_sum[8][26] , \ADDER_IN_from_sum[8][25] , 
        \ADDER_IN_from_sum[8][24] , \ADDER_IN_from_sum[8][23] , 
        \ADDER_IN_from_sum[8][22] , \ADDER_IN_from_sum[8][21] , 
        \ADDER_IN_from_sum[8][20] , \ADDER_IN_from_sum[8][19] , 
        \ADDER_IN_from_sum[8][18] , \ADDER_IN_from_sum[8][17] , 
        \ADDER_IN_from_sum[8][16] , \ADDER_IN_from_sum[8][15] , 
        \ADDER_IN_from_sum[8][14] , \ADDER_IN_from_sum[8][13] , 
        \ADDER_IN_from_sum[8][12] , \ADDER_IN_from_sum[8][11] , 
        \ADDER_IN_from_sum[8][10] , \ADDER_IN_from_sum[8][9] , 
        \ADDER_IN_from_sum[8][8] , \ADDER_IN_from_sum[8][7] , 
        \ADDER_IN_from_sum[8][6] , \ADDER_IN_from_sum[8][5] , 
        \ADDER_IN_from_sum[8][4] , \ADDER_IN_from_sum[8][3] , 
        \ADDER_IN_from_sum[8][2] , \ADDER_IN_from_sum[8][1] , 
        \ADDER_IN_from_sum[8][0] }), .B({\ADDER_IN_from_mux[10][63] , 
        \ADDER_IN_from_mux[10][62] , \ADDER_IN_from_mux[10][61] , 
        \ADDER_IN_from_mux[10][60] , \ADDER_IN_from_mux[10][59] , 
        \ADDER_IN_from_mux[10][58] , \ADDER_IN_from_mux[10][57] , 
        \ADDER_IN_from_mux[10][56] , \ADDER_IN_from_mux[10][55] , 
        \ADDER_IN_from_mux[10][54] , \ADDER_IN_from_mux[10][53] , 
        \ADDER_IN_from_mux[10][52] , \ADDER_IN_from_mux[10][51] , 
        \ADDER_IN_from_mux[10][50] , \ADDER_IN_from_mux[10][49] , 
        \ADDER_IN_from_mux[10][48] , \ADDER_IN_from_mux[10][47] , 
        \ADDER_IN_from_mux[10][46] , \ADDER_IN_from_mux[10][45] , 
        \ADDER_IN_from_mux[10][44] , \ADDER_IN_from_mux[10][43] , 
        \ADDER_IN_from_mux[10][42] , \ADDER_IN_from_mux[10][41] , 
        \ADDER_IN_from_mux[10][40] , \ADDER_IN_from_mux[10][39] , 
        \ADDER_IN_from_mux[10][38] , \ADDER_IN_from_mux[10][37] , 
        \ADDER_IN_from_mux[10][36] , \ADDER_IN_from_mux[10][35] , 
        \ADDER_IN_from_mux[10][34] , \ADDER_IN_from_mux[10][33] , 
        \ADDER_IN_from_mux[10][32] , \ADDER_IN_from_mux[10][31] , 
        \ADDER_IN_from_mux[10][30] , \ADDER_IN_from_mux[10][29] , 
        \ADDER_IN_from_mux[10][28] , \ADDER_IN_from_mux[10][27] , 
        \ADDER_IN_from_mux[10][26] , \ADDER_IN_from_mux[10][25] , 
        \ADDER_IN_from_mux[10][24] , \ADDER_IN_from_mux[10][23] , 
        \ADDER_IN_from_mux[10][22] , \ADDER_IN_from_mux[10][21] , 
        \ADDER_IN_from_mux[10][20] , \ADDER_IN_from_mux[10][19] , 
        \ADDER_IN_from_mux[10][18] , \ADDER_IN_from_mux[10][17] , 
        \ADDER_IN_from_mux[10][16] , \ADDER_IN_from_mux[10][15] , 
        \ADDER_IN_from_mux[10][14] , \ADDER_IN_from_mux[10][13] , 
        \ADDER_IN_from_mux[10][12] , \ADDER_IN_from_mux[10][11] , 
        \ADDER_IN_from_mux[10][10] , \ADDER_IN_from_mux[10][9] , 
        \ADDER_IN_from_mux[10][8] , \ADDER_IN_from_mux[10][7] , 
        \ADDER_IN_from_mux[10][6] , \ADDER_IN_from_mux[10][5] , 
        \ADDER_IN_from_mux[10][4] , \ADDER_IN_from_mux[10][3] , 
        \ADDER_IN_from_mux[10][2] , \ADDER_IN_from_mux[10][1] , 
        \ADDER_IN_from_mux[10][0] }), .S({\ADDER_IN_from_sum[9][63] , 
        \ADDER_IN_from_sum[9][62] , \ADDER_IN_from_sum[9][61] , 
        \ADDER_IN_from_sum[9][60] , \ADDER_IN_from_sum[9][59] , 
        \ADDER_IN_from_sum[9][58] , \ADDER_IN_from_sum[9][57] , 
        \ADDER_IN_from_sum[9][56] , \ADDER_IN_from_sum[9][55] , 
        \ADDER_IN_from_sum[9][54] , \ADDER_IN_from_sum[9][53] , 
        \ADDER_IN_from_sum[9][52] , \ADDER_IN_from_sum[9][51] , 
        \ADDER_IN_from_sum[9][50] , \ADDER_IN_from_sum[9][49] , 
        \ADDER_IN_from_sum[9][48] , \ADDER_IN_from_sum[9][47] , 
        \ADDER_IN_from_sum[9][46] , \ADDER_IN_from_sum[9][45] , 
        \ADDER_IN_from_sum[9][44] , \ADDER_IN_from_sum[9][43] , 
        \ADDER_IN_from_sum[9][42] , \ADDER_IN_from_sum[9][41] , 
        \ADDER_IN_from_sum[9][40] , \ADDER_IN_from_sum[9][39] , 
        \ADDER_IN_from_sum[9][38] , \ADDER_IN_from_sum[9][37] , 
        \ADDER_IN_from_sum[9][36] , \ADDER_IN_from_sum[9][35] , 
        \ADDER_IN_from_sum[9][34] , \ADDER_IN_from_sum[9][33] , 
        \ADDER_IN_from_sum[9][32] , \ADDER_IN_from_sum[9][31] , 
        \ADDER_IN_from_sum[9][30] , \ADDER_IN_from_sum[9][29] , 
        \ADDER_IN_from_sum[9][28] , \ADDER_IN_from_sum[9][27] , 
        \ADDER_IN_from_sum[9][26] , \ADDER_IN_from_sum[9][25] , 
        \ADDER_IN_from_sum[9][24] , \ADDER_IN_from_sum[9][23] , 
        \ADDER_IN_from_sum[9][22] , \ADDER_IN_from_sum[9][21] , 
        \ADDER_IN_from_sum[9][20] , \ADDER_IN_from_sum[9][19] , 
        \ADDER_IN_from_sum[9][18] , \ADDER_IN_from_sum[9][17] , 
        \ADDER_IN_from_sum[9][16] , \ADDER_IN_from_sum[9][15] , 
        \ADDER_IN_from_sum[9][14] , \ADDER_IN_from_sum[9][13] , 
        \ADDER_IN_from_sum[9][12] , \ADDER_IN_from_sum[9][11] , 
        \ADDER_IN_from_sum[9][10] , \ADDER_IN_from_sum[9][9] , 
        \ADDER_IN_from_sum[9][8] , \ADDER_IN_from_sum[9][7] , 
        \ADDER_IN_from_sum[9][6] , \ADDER_IN_from_sum[9][5] , 
        \ADDER_IN_from_sum[9][4] , \ADDER_IN_from_sum[9][3] , 
        \ADDER_IN_from_sum[9][2] , \ADDER_IN_from_sum[9][1] , 
        \ADDER_IN_from_sum[9][0] }) );
  RCA_NBIT64_5 RCA_n_9 ( .A({\ADDER_IN_from_sum[9][63] , 
        \ADDER_IN_from_sum[9][62] , \ADDER_IN_from_sum[9][61] , 
        \ADDER_IN_from_sum[9][60] , \ADDER_IN_from_sum[9][59] , 
        \ADDER_IN_from_sum[9][58] , \ADDER_IN_from_sum[9][57] , 
        \ADDER_IN_from_sum[9][56] , \ADDER_IN_from_sum[9][55] , 
        \ADDER_IN_from_sum[9][54] , \ADDER_IN_from_sum[9][53] , 
        \ADDER_IN_from_sum[9][52] , \ADDER_IN_from_sum[9][51] , 
        \ADDER_IN_from_sum[9][50] , \ADDER_IN_from_sum[9][49] , 
        \ADDER_IN_from_sum[9][48] , \ADDER_IN_from_sum[9][47] , 
        \ADDER_IN_from_sum[9][46] , \ADDER_IN_from_sum[9][45] , 
        \ADDER_IN_from_sum[9][44] , \ADDER_IN_from_sum[9][43] , 
        \ADDER_IN_from_sum[9][42] , \ADDER_IN_from_sum[9][41] , 
        \ADDER_IN_from_sum[9][40] , \ADDER_IN_from_sum[9][39] , 
        \ADDER_IN_from_sum[9][38] , \ADDER_IN_from_sum[9][37] , 
        \ADDER_IN_from_sum[9][36] , \ADDER_IN_from_sum[9][35] , 
        \ADDER_IN_from_sum[9][34] , \ADDER_IN_from_sum[9][33] , 
        \ADDER_IN_from_sum[9][32] , \ADDER_IN_from_sum[9][31] , 
        \ADDER_IN_from_sum[9][30] , \ADDER_IN_from_sum[9][29] , 
        \ADDER_IN_from_sum[9][28] , \ADDER_IN_from_sum[9][27] , 
        \ADDER_IN_from_sum[9][26] , \ADDER_IN_from_sum[9][25] , 
        \ADDER_IN_from_sum[9][24] , \ADDER_IN_from_sum[9][23] , 
        \ADDER_IN_from_sum[9][22] , \ADDER_IN_from_sum[9][21] , 
        \ADDER_IN_from_sum[9][20] , \ADDER_IN_from_sum[9][19] , 
        \ADDER_IN_from_sum[9][18] , \ADDER_IN_from_sum[9][17] , 
        \ADDER_IN_from_sum[9][16] , \ADDER_IN_from_sum[9][15] , 
        \ADDER_IN_from_sum[9][14] , \ADDER_IN_from_sum[9][13] , 
        \ADDER_IN_from_sum[9][12] , \ADDER_IN_from_sum[9][11] , 
        \ADDER_IN_from_sum[9][10] , \ADDER_IN_from_sum[9][9] , 
        \ADDER_IN_from_sum[9][8] , \ADDER_IN_from_sum[9][7] , 
        \ADDER_IN_from_sum[9][6] , \ADDER_IN_from_sum[9][5] , 
        \ADDER_IN_from_sum[9][4] , \ADDER_IN_from_sum[9][3] , 
        \ADDER_IN_from_sum[9][2] , \ADDER_IN_from_sum[9][1] , 
        \ADDER_IN_from_sum[9][0] }), .B({\ADDER_IN_from_mux[11][63] , 
        \ADDER_IN_from_mux[11][62] , \ADDER_IN_from_mux[11][61] , 
        \ADDER_IN_from_mux[11][60] , \ADDER_IN_from_mux[11][59] , 
        \ADDER_IN_from_mux[11][58] , \ADDER_IN_from_mux[11][57] , 
        \ADDER_IN_from_mux[11][56] , \ADDER_IN_from_mux[11][55] , 
        \ADDER_IN_from_mux[11][54] , \ADDER_IN_from_mux[11][53] , 
        \ADDER_IN_from_mux[11][52] , \ADDER_IN_from_mux[11][51] , 
        \ADDER_IN_from_mux[11][50] , \ADDER_IN_from_mux[11][49] , 
        \ADDER_IN_from_mux[11][48] , \ADDER_IN_from_mux[11][47] , 
        \ADDER_IN_from_mux[11][46] , \ADDER_IN_from_mux[11][45] , 
        \ADDER_IN_from_mux[11][44] , \ADDER_IN_from_mux[11][43] , 
        \ADDER_IN_from_mux[11][42] , \ADDER_IN_from_mux[11][41] , 
        \ADDER_IN_from_mux[11][40] , \ADDER_IN_from_mux[11][39] , 
        \ADDER_IN_from_mux[11][38] , \ADDER_IN_from_mux[11][37] , 
        \ADDER_IN_from_mux[11][36] , \ADDER_IN_from_mux[11][35] , 
        \ADDER_IN_from_mux[11][34] , \ADDER_IN_from_mux[11][33] , 
        \ADDER_IN_from_mux[11][32] , \ADDER_IN_from_mux[11][31] , 
        \ADDER_IN_from_mux[11][30] , \ADDER_IN_from_mux[11][29] , 
        \ADDER_IN_from_mux[11][28] , \ADDER_IN_from_mux[11][27] , 
        \ADDER_IN_from_mux[11][26] , \ADDER_IN_from_mux[11][25] , 
        \ADDER_IN_from_mux[11][24] , \ADDER_IN_from_mux[11][23] , 
        \ADDER_IN_from_mux[11][22] , \ADDER_IN_from_mux[11][21] , 
        \ADDER_IN_from_mux[11][20] , \ADDER_IN_from_mux[11][19] , 
        \ADDER_IN_from_mux[11][18] , \ADDER_IN_from_mux[11][17] , 
        \ADDER_IN_from_mux[11][16] , \ADDER_IN_from_mux[11][15] , 
        \ADDER_IN_from_mux[11][14] , \ADDER_IN_from_mux[11][13] , 
        \ADDER_IN_from_mux[11][12] , \ADDER_IN_from_mux[11][11] , 
        \ADDER_IN_from_mux[11][10] , \ADDER_IN_from_mux[11][9] , 
        \ADDER_IN_from_mux[11][8] , \ADDER_IN_from_mux[11][7] , 
        \ADDER_IN_from_mux[11][6] , \ADDER_IN_from_mux[11][5] , 
        \ADDER_IN_from_mux[11][4] , \ADDER_IN_from_mux[11][3] , 
        \ADDER_IN_from_mux[11][2] , \ADDER_IN_from_mux[11][1] , 
        \ADDER_IN_from_mux[11][0] }), .S({\ADDER_IN_from_sum[10][63] , 
        \ADDER_IN_from_sum[10][62] , \ADDER_IN_from_sum[10][61] , 
        \ADDER_IN_from_sum[10][60] , \ADDER_IN_from_sum[10][59] , 
        \ADDER_IN_from_sum[10][58] , \ADDER_IN_from_sum[10][57] , 
        \ADDER_IN_from_sum[10][56] , \ADDER_IN_from_sum[10][55] , 
        \ADDER_IN_from_sum[10][54] , \ADDER_IN_from_sum[10][53] , 
        \ADDER_IN_from_sum[10][52] , \ADDER_IN_from_sum[10][51] , 
        \ADDER_IN_from_sum[10][50] , \ADDER_IN_from_sum[10][49] , 
        \ADDER_IN_from_sum[10][48] , \ADDER_IN_from_sum[10][47] , 
        \ADDER_IN_from_sum[10][46] , \ADDER_IN_from_sum[10][45] , 
        \ADDER_IN_from_sum[10][44] , \ADDER_IN_from_sum[10][43] , 
        \ADDER_IN_from_sum[10][42] , \ADDER_IN_from_sum[10][41] , 
        \ADDER_IN_from_sum[10][40] , \ADDER_IN_from_sum[10][39] , 
        \ADDER_IN_from_sum[10][38] , \ADDER_IN_from_sum[10][37] , 
        \ADDER_IN_from_sum[10][36] , \ADDER_IN_from_sum[10][35] , 
        \ADDER_IN_from_sum[10][34] , \ADDER_IN_from_sum[10][33] , 
        \ADDER_IN_from_sum[10][32] , \ADDER_IN_from_sum[10][31] , 
        \ADDER_IN_from_sum[10][30] , \ADDER_IN_from_sum[10][29] , 
        \ADDER_IN_from_sum[10][28] , \ADDER_IN_from_sum[10][27] , 
        \ADDER_IN_from_sum[10][26] , \ADDER_IN_from_sum[10][25] , 
        \ADDER_IN_from_sum[10][24] , \ADDER_IN_from_sum[10][23] , 
        \ADDER_IN_from_sum[10][22] , \ADDER_IN_from_sum[10][21] , 
        \ADDER_IN_from_sum[10][20] , \ADDER_IN_from_sum[10][19] , 
        \ADDER_IN_from_sum[10][18] , \ADDER_IN_from_sum[10][17] , 
        \ADDER_IN_from_sum[10][16] , \ADDER_IN_from_sum[10][15] , 
        \ADDER_IN_from_sum[10][14] , \ADDER_IN_from_sum[10][13] , 
        \ADDER_IN_from_sum[10][12] , \ADDER_IN_from_sum[10][11] , 
        \ADDER_IN_from_sum[10][10] , \ADDER_IN_from_sum[10][9] , 
        \ADDER_IN_from_sum[10][8] , \ADDER_IN_from_sum[10][7] , 
        \ADDER_IN_from_sum[10][6] , \ADDER_IN_from_sum[10][5] , 
        \ADDER_IN_from_sum[10][4] , \ADDER_IN_from_sum[10][3] , 
        \ADDER_IN_from_sum[10][2] , \ADDER_IN_from_sum[10][1] , 
        \ADDER_IN_from_sum[10][0] }) );
  RCA_NBIT64_4 RCA_n_10 ( .A({\ADDER_IN_from_sum[10][63] , 
        \ADDER_IN_from_sum[10][62] , \ADDER_IN_from_sum[10][61] , 
        \ADDER_IN_from_sum[10][60] , \ADDER_IN_from_sum[10][59] , 
        \ADDER_IN_from_sum[10][58] , \ADDER_IN_from_sum[10][57] , 
        \ADDER_IN_from_sum[10][56] , \ADDER_IN_from_sum[10][55] , 
        \ADDER_IN_from_sum[10][54] , \ADDER_IN_from_sum[10][53] , 
        \ADDER_IN_from_sum[10][52] , \ADDER_IN_from_sum[10][51] , 
        \ADDER_IN_from_sum[10][50] , \ADDER_IN_from_sum[10][49] , 
        \ADDER_IN_from_sum[10][48] , \ADDER_IN_from_sum[10][47] , 
        \ADDER_IN_from_sum[10][46] , \ADDER_IN_from_sum[10][45] , 
        \ADDER_IN_from_sum[10][44] , \ADDER_IN_from_sum[10][43] , 
        \ADDER_IN_from_sum[10][42] , \ADDER_IN_from_sum[10][41] , 
        \ADDER_IN_from_sum[10][40] , \ADDER_IN_from_sum[10][39] , 
        \ADDER_IN_from_sum[10][38] , \ADDER_IN_from_sum[10][37] , 
        \ADDER_IN_from_sum[10][36] , \ADDER_IN_from_sum[10][35] , 
        \ADDER_IN_from_sum[10][34] , \ADDER_IN_from_sum[10][33] , 
        \ADDER_IN_from_sum[10][32] , \ADDER_IN_from_sum[10][31] , 
        \ADDER_IN_from_sum[10][30] , \ADDER_IN_from_sum[10][29] , 
        \ADDER_IN_from_sum[10][28] , \ADDER_IN_from_sum[10][27] , 
        \ADDER_IN_from_sum[10][26] , \ADDER_IN_from_sum[10][25] , 
        \ADDER_IN_from_sum[10][24] , \ADDER_IN_from_sum[10][23] , 
        \ADDER_IN_from_sum[10][22] , \ADDER_IN_from_sum[10][21] , 
        \ADDER_IN_from_sum[10][20] , \ADDER_IN_from_sum[10][19] , 
        \ADDER_IN_from_sum[10][18] , \ADDER_IN_from_sum[10][17] , 
        \ADDER_IN_from_sum[10][16] , \ADDER_IN_from_sum[10][15] , 
        \ADDER_IN_from_sum[10][14] , \ADDER_IN_from_sum[10][13] , 
        \ADDER_IN_from_sum[10][12] , \ADDER_IN_from_sum[10][11] , 
        \ADDER_IN_from_sum[10][10] , \ADDER_IN_from_sum[10][9] , 
        \ADDER_IN_from_sum[10][8] , \ADDER_IN_from_sum[10][7] , 
        \ADDER_IN_from_sum[10][6] , \ADDER_IN_from_sum[10][5] , 
        \ADDER_IN_from_sum[10][4] , \ADDER_IN_from_sum[10][3] , 
        \ADDER_IN_from_sum[10][2] , \ADDER_IN_from_sum[10][1] , 
        \ADDER_IN_from_sum[10][0] }), .B({\ADDER_IN_from_mux[12][63] , 
        \ADDER_IN_from_mux[12][62] , \ADDER_IN_from_mux[12][61] , 
        \ADDER_IN_from_mux[12][60] , \ADDER_IN_from_mux[12][59] , 
        \ADDER_IN_from_mux[12][58] , \ADDER_IN_from_mux[12][57] , 
        \ADDER_IN_from_mux[12][56] , \ADDER_IN_from_mux[12][55] , 
        \ADDER_IN_from_mux[12][54] , \ADDER_IN_from_mux[12][53] , 
        \ADDER_IN_from_mux[12][52] , \ADDER_IN_from_mux[12][51] , 
        \ADDER_IN_from_mux[12][50] , \ADDER_IN_from_mux[12][49] , 
        \ADDER_IN_from_mux[12][48] , \ADDER_IN_from_mux[12][47] , 
        \ADDER_IN_from_mux[12][46] , \ADDER_IN_from_mux[12][45] , 
        \ADDER_IN_from_mux[12][44] , \ADDER_IN_from_mux[12][43] , 
        \ADDER_IN_from_mux[12][42] , \ADDER_IN_from_mux[12][41] , 
        \ADDER_IN_from_mux[12][40] , \ADDER_IN_from_mux[12][39] , 
        \ADDER_IN_from_mux[12][38] , \ADDER_IN_from_mux[12][37] , 
        \ADDER_IN_from_mux[12][36] , \ADDER_IN_from_mux[12][35] , 
        \ADDER_IN_from_mux[12][34] , \ADDER_IN_from_mux[12][33] , 
        \ADDER_IN_from_mux[12][32] , \ADDER_IN_from_mux[12][31] , 
        \ADDER_IN_from_mux[12][30] , \ADDER_IN_from_mux[12][29] , 
        \ADDER_IN_from_mux[12][28] , \ADDER_IN_from_mux[12][27] , 
        \ADDER_IN_from_mux[12][26] , \ADDER_IN_from_mux[12][25] , 
        \ADDER_IN_from_mux[12][24] , \ADDER_IN_from_mux[12][23] , 
        \ADDER_IN_from_mux[12][22] , \ADDER_IN_from_mux[12][21] , 
        \ADDER_IN_from_mux[12][20] , \ADDER_IN_from_mux[12][19] , 
        \ADDER_IN_from_mux[12][18] , \ADDER_IN_from_mux[12][17] , 
        \ADDER_IN_from_mux[12][16] , \ADDER_IN_from_mux[12][15] , 
        \ADDER_IN_from_mux[12][14] , \ADDER_IN_from_mux[12][13] , 
        \ADDER_IN_from_mux[12][12] , \ADDER_IN_from_mux[12][11] , 
        \ADDER_IN_from_mux[12][10] , \ADDER_IN_from_mux[12][9] , 
        \ADDER_IN_from_mux[12][8] , \ADDER_IN_from_mux[12][7] , 
        \ADDER_IN_from_mux[12][6] , \ADDER_IN_from_mux[12][5] , 
        \ADDER_IN_from_mux[12][4] , \ADDER_IN_from_mux[12][3] , 
        \ADDER_IN_from_mux[12][2] , \ADDER_IN_from_mux[12][1] , 
        \ADDER_IN_from_mux[12][0] }), .S({\ADDER_IN_from_sum[11][63] , 
        \ADDER_IN_from_sum[11][62] , \ADDER_IN_from_sum[11][61] , 
        \ADDER_IN_from_sum[11][60] , \ADDER_IN_from_sum[11][59] , 
        \ADDER_IN_from_sum[11][58] , \ADDER_IN_from_sum[11][57] , 
        \ADDER_IN_from_sum[11][56] , \ADDER_IN_from_sum[11][55] , 
        \ADDER_IN_from_sum[11][54] , \ADDER_IN_from_sum[11][53] , 
        \ADDER_IN_from_sum[11][52] , \ADDER_IN_from_sum[11][51] , 
        \ADDER_IN_from_sum[11][50] , \ADDER_IN_from_sum[11][49] , 
        \ADDER_IN_from_sum[11][48] , \ADDER_IN_from_sum[11][47] , 
        \ADDER_IN_from_sum[11][46] , \ADDER_IN_from_sum[11][45] , 
        \ADDER_IN_from_sum[11][44] , \ADDER_IN_from_sum[11][43] , 
        \ADDER_IN_from_sum[11][42] , \ADDER_IN_from_sum[11][41] , 
        \ADDER_IN_from_sum[11][40] , \ADDER_IN_from_sum[11][39] , 
        \ADDER_IN_from_sum[11][38] , \ADDER_IN_from_sum[11][37] , 
        \ADDER_IN_from_sum[11][36] , \ADDER_IN_from_sum[11][35] , 
        \ADDER_IN_from_sum[11][34] , \ADDER_IN_from_sum[11][33] , 
        \ADDER_IN_from_sum[11][32] , \ADDER_IN_from_sum[11][31] , 
        \ADDER_IN_from_sum[11][30] , \ADDER_IN_from_sum[11][29] , 
        \ADDER_IN_from_sum[11][28] , \ADDER_IN_from_sum[11][27] , 
        \ADDER_IN_from_sum[11][26] , \ADDER_IN_from_sum[11][25] , 
        \ADDER_IN_from_sum[11][24] , \ADDER_IN_from_sum[11][23] , 
        \ADDER_IN_from_sum[11][22] , \ADDER_IN_from_sum[11][21] , 
        \ADDER_IN_from_sum[11][20] , \ADDER_IN_from_sum[11][19] , 
        \ADDER_IN_from_sum[11][18] , \ADDER_IN_from_sum[11][17] , 
        \ADDER_IN_from_sum[11][16] , \ADDER_IN_from_sum[11][15] , 
        \ADDER_IN_from_sum[11][14] , \ADDER_IN_from_sum[11][13] , 
        \ADDER_IN_from_sum[11][12] , \ADDER_IN_from_sum[11][11] , 
        \ADDER_IN_from_sum[11][10] , \ADDER_IN_from_sum[11][9] , 
        \ADDER_IN_from_sum[11][8] , \ADDER_IN_from_sum[11][7] , 
        \ADDER_IN_from_sum[11][6] , \ADDER_IN_from_sum[11][5] , 
        \ADDER_IN_from_sum[11][4] , \ADDER_IN_from_sum[11][3] , 
        \ADDER_IN_from_sum[11][2] , \ADDER_IN_from_sum[11][1] , 
        \ADDER_IN_from_sum[11][0] }) );
  RCA_NBIT64_3 RCA_n_11 ( .A({\ADDER_IN_from_sum[11][63] , 
        \ADDER_IN_from_sum[11][62] , \ADDER_IN_from_sum[11][61] , 
        \ADDER_IN_from_sum[11][60] , \ADDER_IN_from_sum[11][59] , 
        \ADDER_IN_from_sum[11][58] , \ADDER_IN_from_sum[11][57] , 
        \ADDER_IN_from_sum[11][56] , \ADDER_IN_from_sum[11][55] , 
        \ADDER_IN_from_sum[11][54] , \ADDER_IN_from_sum[11][53] , 
        \ADDER_IN_from_sum[11][52] , \ADDER_IN_from_sum[11][51] , 
        \ADDER_IN_from_sum[11][50] , \ADDER_IN_from_sum[11][49] , 
        \ADDER_IN_from_sum[11][48] , \ADDER_IN_from_sum[11][47] , 
        \ADDER_IN_from_sum[11][46] , \ADDER_IN_from_sum[11][45] , 
        \ADDER_IN_from_sum[11][44] , \ADDER_IN_from_sum[11][43] , 
        \ADDER_IN_from_sum[11][42] , \ADDER_IN_from_sum[11][41] , 
        \ADDER_IN_from_sum[11][40] , \ADDER_IN_from_sum[11][39] , 
        \ADDER_IN_from_sum[11][38] , \ADDER_IN_from_sum[11][37] , 
        \ADDER_IN_from_sum[11][36] , \ADDER_IN_from_sum[11][35] , 
        \ADDER_IN_from_sum[11][34] , \ADDER_IN_from_sum[11][33] , 
        \ADDER_IN_from_sum[11][32] , \ADDER_IN_from_sum[11][31] , 
        \ADDER_IN_from_sum[11][30] , \ADDER_IN_from_sum[11][29] , 
        \ADDER_IN_from_sum[11][28] , \ADDER_IN_from_sum[11][27] , 
        \ADDER_IN_from_sum[11][26] , \ADDER_IN_from_sum[11][25] , 
        \ADDER_IN_from_sum[11][24] , \ADDER_IN_from_sum[11][23] , 
        \ADDER_IN_from_sum[11][22] , \ADDER_IN_from_sum[11][21] , 
        \ADDER_IN_from_sum[11][20] , \ADDER_IN_from_sum[11][19] , 
        \ADDER_IN_from_sum[11][18] , \ADDER_IN_from_sum[11][17] , 
        \ADDER_IN_from_sum[11][16] , \ADDER_IN_from_sum[11][15] , 
        \ADDER_IN_from_sum[11][14] , \ADDER_IN_from_sum[11][13] , 
        \ADDER_IN_from_sum[11][12] , \ADDER_IN_from_sum[11][11] , 
        \ADDER_IN_from_sum[11][10] , \ADDER_IN_from_sum[11][9] , 
        \ADDER_IN_from_sum[11][8] , \ADDER_IN_from_sum[11][7] , 
        \ADDER_IN_from_sum[11][6] , \ADDER_IN_from_sum[11][5] , 
        \ADDER_IN_from_sum[11][4] , \ADDER_IN_from_sum[11][3] , 
        \ADDER_IN_from_sum[11][2] , \ADDER_IN_from_sum[11][1] , 
        \ADDER_IN_from_sum[11][0] }), .B({\ADDER_IN_from_mux[13][63] , 
        \ADDER_IN_from_mux[13][62] , \ADDER_IN_from_mux[13][61] , 
        \ADDER_IN_from_mux[13][60] , \ADDER_IN_from_mux[13][59] , 
        \ADDER_IN_from_mux[13][58] , \ADDER_IN_from_mux[13][57] , 
        \ADDER_IN_from_mux[13][56] , \ADDER_IN_from_mux[13][55] , 
        \ADDER_IN_from_mux[13][54] , \ADDER_IN_from_mux[13][53] , 
        \ADDER_IN_from_mux[13][52] , \ADDER_IN_from_mux[13][51] , 
        \ADDER_IN_from_mux[13][50] , \ADDER_IN_from_mux[13][49] , 
        \ADDER_IN_from_mux[13][48] , \ADDER_IN_from_mux[13][47] , 
        \ADDER_IN_from_mux[13][46] , \ADDER_IN_from_mux[13][45] , 
        \ADDER_IN_from_mux[13][44] , \ADDER_IN_from_mux[13][43] , 
        \ADDER_IN_from_mux[13][42] , \ADDER_IN_from_mux[13][41] , 
        \ADDER_IN_from_mux[13][40] , \ADDER_IN_from_mux[13][39] , 
        \ADDER_IN_from_mux[13][38] , \ADDER_IN_from_mux[13][37] , 
        \ADDER_IN_from_mux[13][36] , \ADDER_IN_from_mux[13][35] , 
        \ADDER_IN_from_mux[13][34] , \ADDER_IN_from_mux[13][33] , 
        \ADDER_IN_from_mux[13][32] , \ADDER_IN_from_mux[13][31] , 
        \ADDER_IN_from_mux[13][30] , \ADDER_IN_from_mux[13][29] , 
        \ADDER_IN_from_mux[13][28] , \ADDER_IN_from_mux[13][27] , 
        \ADDER_IN_from_mux[13][26] , \ADDER_IN_from_mux[13][25] , 
        \ADDER_IN_from_mux[13][24] , \ADDER_IN_from_mux[13][23] , 
        \ADDER_IN_from_mux[13][22] , \ADDER_IN_from_mux[13][21] , 
        \ADDER_IN_from_mux[13][20] , \ADDER_IN_from_mux[13][19] , 
        \ADDER_IN_from_mux[13][18] , \ADDER_IN_from_mux[13][17] , 
        \ADDER_IN_from_mux[13][16] , \ADDER_IN_from_mux[13][15] , 
        \ADDER_IN_from_mux[13][14] , \ADDER_IN_from_mux[13][13] , 
        \ADDER_IN_from_mux[13][12] , \ADDER_IN_from_mux[13][11] , 
        \ADDER_IN_from_mux[13][10] , \ADDER_IN_from_mux[13][9] , 
        \ADDER_IN_from_mux[13][8] , \ADDER_IN_from_mux[13][7] , 
        \ADDER_IN_from_mux[13][6] , \ADDER_IN_from_mux[13][5] , 
        \ADDER_IN_from_mux[13][4] , \ADDER_IN_from_mux[13][3] , 
        \ADDER_IN_from_mux[13][2] , \ADDER_IN_from_mux[13][1] , 
        \ADDER_IN_from_mux[13][0] }), .S({\ADDER_IN_from_sum[12][63] , 
        \ADDER_IN_from_sum[12][62] , \ADDER_IN_from_sum[12][61] , 
        \ADDER_IN_from_sum[12][60] , \ADDER_IN_from_sum[12][59] , 
        \ADDER_IN_from_sum[12][58] , \ADDER_IN_from_sum[12][57] , 
        \ADDER_IN_from_sum[12][56] , \ADDER_IN_from_sum[12][55] , 
        \ADDER_IN_from_sum[12][54] , \ADDER_IN_from_sum[12][53] , 
        \ADDER_IN_from_sum[12][52] , \ADDER_IN_from_sum[12][51] , 
        \ADDER_IN_from_sum[12][50] , \ADDER_IN_from_sum[12][49] , 
        \ADDER_IN_from_sum[12][48] , \ADDER_IN_from_sum[12][47] , 
        \ADDER_IN_from_sum[12][46] , \ADDER_IN_from_sum[12][45] , 
        \ADDER_IN_from_sum[12][44] , \ADDER_IN_from_sum[12][43] , 
        \ADDER_IN_from_sum[12][42] , \ADDER_IN_from_sum[12][41] , 
        \ADDER_IN_from_sum[12][40] , \ADDER_IN_from_sum[12][39] , 
        \ADDER_IN_from_sum[12][38] , \ADDER_IN_from_sum[12][37] , 
        \ADDER_IN_from_sum[12][36] , \ADDER_IN_from_sum[12][35] , 
        \ADDER_IN_from_sum[12][34] , \ADDER_IN_from_sum[12][33] , 
        \ADDER_IN_from_sum[12][32] , \ADDER_IN_from_sum[12][31] , 
        \ADDER_IN_from_sum[12][30] , \ADDER_IN_from_sum[12][29] , 
        \ADDER_IN_from_sum[12][28] , \ADDER_IN_from_sum[12][27] , 
        \ADDER_IN_from_sum[12][26] , \ADDER_IN_from_sum[12][25] , 
        \ADDER_IN_from_sum[12][24] , \ADDER_IN_from_sum[12][23] , 
        \ADDER_IN_from_sum[12][22] , \ADDER_IN_from_sum[12][21] , 
        \ADDER_IN_from_sum[12][20] , \ADDER_IN_from_sum[12][19] , 
        \ADDER_IN_from_sum[12][18] , \ADDER_IN_from_sum[12][17] , 
        \ADDER_IN_from_sum[12][16] , \ADDER_IN_from_sum[12][15] , 
        \ADDER_IN_from_sum[12][14] , \ADDER_IN_from_sum[12][13] , 
        \ADDER_IN_from_sum[12][12] , \ADDER_IN_from_sum[12][11] , 
        \ADDER_IN_from_sum[12][10] , \ADDER_IN_from_sum[12][9] , 
        \ADDER_IN_from_sum[12][8] , \ADDER_IN_from_sum[12][7] , 
        \ADDER_IN_from_sum[12][6] , \ADDER_IN_from_sum[12][5] , 
        \ADDER_IN_from_sum[12][4] , \ADDER_IN_from_sum[12][3] , 
        \ADDER_IN_from_sum[12][2] , \ADDER_IN_from_sum[12][1] , 
        \ADDER_IN_from_sum[12][0] }) );
  RCA_NBIT64_2 RCA_n_12 ( .A({\ADDER_IN_from_sum[12][63] , 
        \ADDER_IN_from_sum[12][62] , \ADDER_IN_from_sum[12][61] , 
        \ADDER_IN_from_sum[12][60] , \ADDER_IN_from_sum[12][59] , 
        \ADDER_IN_from_sum[12][58] , \ADDER_IN_from_sum[12][57] , 
        \ADDER_IN_from_sum[12][56] , \ADDER_IN_from_sum[12][55] , 
        \ADDER_IN_from_sum[12][54] , \ADDER_IN_from_sum[12][53] , 
        \ADDER_IN_from_sum[12][52] , \ADDER_IN_from_sum[12][51] , 
        \ADDER_IN_from_sum[12][50] , \ADDER_IN_from_sum[12][49] , 
        \ADDER_IN_from_sum[12][48] , \ADDER_IN_from_sum[12][47] , 
        \ADDER_IN_from_sum[12][46] , \ADDER_IN_from_sum[12][45] , 
        \ADDER_IN_from_sum[12][44] , \ADDER_IN_from_sum[12][43] , 
        \ADDER_IN_from_sum[12][42] , \ADDER_IN_from_sum[12][41] , 
        \ADDER_IN_from_sum[12][40] , \ADDER_IN_from_sum[12][39] , 
        \ADDER_IN_from_sum[12][38] , \ADDER_IN_from_sum[12][37] , 
        \ADDER_IN_from_sum[12][36] , \ADDER_IN_from_sum[12][35] , 
        \ADDER_IN_from_sum[12][34] , \ADDER_IN_from_sum[12][33] , 
        \ADDER_IN_from_sum[12][32] , \ADDER_IN_from_sum[12][31] , 
        \ADDER_IN_from_sum[12][30] , \ADDER_IN_from_sum[12][29] , 
        \ADDER_IN_from_sum[12][28] , \ADDER_IN_from_sum[12][27] , 
        \ADDER_IN_from_sum[12][26] , \ADDER_IN_from_sum[12][25] , 
        \ADDER_IN_from_sum[12][24] , \ADDER_IN_from_sum[12][23] , 
        \ADDER_IN_from_sum[12][22] , \ADDER_IN_from_sum[12][21] , 
        \ADDER_IN_from_sum[12][20] , \ADDER_IN_from_sum[12][19] , 
        \ADDER_IN_from_sum[12][18] , \ADDER_IN_from_sum[12][17] , 
        \ADDER_IN_from_sum[12][16] , \ADDER_IN_from_sum[12][15] , 
        \ADDER_IN_from_sum[12][14] , \ADDER_IN_from_sum[12][13] , 
        \ADDER_IN_from_sum[12][12] , \ADDER_IN_from_sum[12][11] , 
        \ADDER_IN_from_sum[12][10] , \ADDER_IN_from_sum[12][9] , 
        \ADDER_IN_from_sum[12][8] , \ADDER_IN_from_sum[12][7] , 
        \ADDER_IN_from_sum[12][6] , \ADDER_IN_from_sum[12][5] , 
        \ADDER_IN_from_sum[12][4] , \ADDER_IN_from_sum[12][3] , 
        \ADDER_IN_from_sum[12][2] , \ADDER_IN_from_sum[12][1] , 
        \ADDER_IN_from_sum[12][0] }), .B({\ADDER_IN_from_mux[14][63] , 
        \ADDER_IN_from_mux[14][62] , \ADDER_IN_from_mux[14][61] , 
        \ADDER_IN_from_mux[14][60] , \ADDER_IN_from_mux[14][59] , 
        \ADDER_IN_from_mux[14][58] , \ADDER_IN_from_mux[14][57] , 
        \ADDER_IN_from_mux[14][56] , \ADDER_IN_from_mux[14][55] , 
        \ADDER_IN_from_mux[14][54] , \ADDER_IN_from_mux[14][53] , 
        \ADDER_IN_from_mux[14][52] , \ADDER_IN_from_mux[14][51] , 
        \ADDER_IN_from_mux[14][50] , \ADDER_IN_from_mux[14][49] , 
        \ADDER_IN_from_mux[14][48] , \ADDER_IN_from_mux[14][47] , 
        \ADDER_IN_from_mux[14][46] , \ADDER_IN_from_mux[14][45] , 
        \ADDER_IN_from_mux[14][44] , \ADDER_IN_from_mux[14][43] , 
        \ADDER_IN_from_mux[14][42] , \ADDER_IN_from_mux[14][41] , 
        \ADDER_IN_from_mux[14][40] , \ADDER_IN_from_mux[14][39] , 
        \ADDER_IN_from_mux[14][38] , \ADDER_IN_from_mux[14][37] , 
        \ADDER_IN_from_mux[14][36] , \ADDER_IN_from_mux[14][35] , 
        \ADDER_IN_from_mux[14][34] , \ADDER_IN_from_mux[14][33] , 
        \ADDER_IN_from_mux[14][32] , \ADDER_IN_from_mux[14][31] , 
        \ADDER_IN_from_mux[14][30] , \ADDER_IN_from_mux[14][29] , 
        \ADDER_IN_from_mux[14][28] , \ADDER_IN_from_mux[14][27] , 
        \ADDER_IN_from_mux[14][26] , \ADDER_IN_from_mux[14][25] , 
        \ADDER_IN_from_mux[14][24] , \ADDER_IN_from_mux[14][23] , 
        \ADDER_IN_from_mux[14][22] , \ADDER_IN_from_mux[14][21] , 
        \ADDER_IN_from_mux[14][20] , \ADDER_IN_from_mux[14][19] , 
        \ADDER_IN_from_mux[14][18] , \ADDER_IN_from_mux[14][17] , 
        \ADDER_IN_from_mux[14][16] , \ADDER_IN_from_mux[14][15] , 
        \ADDER_IN_from_mux[14][14] , \ADDER_IN_from_mux[14][13] , 
        \ADDER_IN_from_mux[14][12] , \ADDER_IN_from_mux[14][11] , 
        \ADDER_IN_from_mux[14][10] , \ADDER_IN_from_mux[14][9] , 
        \ADDER_IN_from_mux[14][8] , \ADDER_IN_from_mux[14][7] , 
        \ADDER_IN_from_mux[14][6] , \ADDER_IN_from_mux[14][5] , 
        \ADDER_IN_from_mux[14][4] , \ADDER_IN_from_mux[14][3] , 
        \ADDER_IN_from_mux[14][2] , \ADDER_IN_from_mux[14][1] , 
        \ADDER_IN_from_mux[14][0] }), .S({\ADDER_IN_from_sum[13][63] , 
        \ADDER_IN_from_sum[13][62] , \ADDER_IN_from_sum[13][61] , 
        \ADDER_IN_from_sum[13][60] , \ADDER_IN_from_sum[13][59] , 
        \ADDER_IN_from_sum[13][58] , \ADDER_IN_from_sum[13][57] , 
        \ADDER_IN_from_sum[13][56] , \ADDER_IN_from_sum[13][55] , 
        \ADDER_IN_from_sum[13][54] , \ADDER_IN_from_sum[13][53] , 
        \ADDER_IN_from_sum[13][52] , \ADDER_IN_from_sum[13][51] , 
        \ADDER_IN_from_sum[13][50] , \ADDER_IN_from_sum[13][49] , 
        \ADDER_IN_from_sum[13][48] , \ADDER_IN_from_sum[13][47] , 
        \ADDER_IN_from_sum[13][46] , \ADDER_IN_from_sum[13][45] , 
        \ADDER_IN_from_sum[13][44] , \ADDER_IN_from_sum[13][43] , 
        \ADDER_IN_from_sum[13][42] , \ADDER_IN_from_sum[13][41] , 
        \ADDER_IN_from_sum[13][40] , \ADDER_IN_from_sum[13][39] , 
        \ADDER_IN_from_sum[13][38] , \ADDER_IN_from_sum[13][37] , 
        \ADDER_IN_from_sum[13][36] , \ADDER_IN_from_sum[13][35] , 
        \ADDER_IN_from_sum[13][34] , \ADDER_IN_from_sum[13][33] , 
        \ADDER_IN_from_sum[13][32] , \ADDER_IN_from_sum[13][31] , 
        \ADDER_IN_from_sum[13][30] , \ADDER_IN_from_sum[13][29] , 
        \ADDER_IN_from_sum[13][28] , \ADDER_IN_from_sum[13][27] , 
        \ADDER_IN_from_sum[13][26] , \ADDER_IN_from_sum[13][25] , 
        \ADDER_IN_from_sum[13][24] , \ADDER_IN_from_sum[13][23] , 
        \ADDER_IN_from_sum[13][22] , \ADDER_IN_from_sum[13][21] , 
        \ADDER_IN_from_sum[13][20] , \ADDER_IN_from_sum[13][19] , 
        \ADDER_IN_from_sum[13][18] , \ADDER_IN_from_sum[13][17] , 
        \ADDER_IN_from_sum[13][16] , \ADDER_IN_from_sum[13][15] , 
        \ADDER_IN_from_sum[13][14] , \ADDER_IN_from_sum[13][13] , 
        \ADDER_IN_from_sum[13][12] , \ADDER_IN_from_sum[13][11] , 
        \ADDER_IN_from_sum[13][10] , \ADDER_IN_from_sum[13][9] , 
        \ADDER_IN_from_sum[13][8] , \ADDER_IN_from_sum[13][7] , 
        \ADDER_IN_from_sum[13][6] , \ADDER_IN_from_sum[13][5] , 
        \ADDER_IN_from_sum[13][4] , \ADDER_IN_from_sum[13][3] , 
        \ADDER_IN_from_sum[13][2] , \ADDER_IN_from_sum[13][1] , 
        \ADDER_IN_from_sum[13][0] }) );
  RCA_NBIT64_1 RCA_n_13 ( .A({\ADDER_IN_from_sum[13][63] , 
        \ADDER_IN_from_sum[13][62] , \ADDER_IN_from_sum[13][61] , 
        \ADDER_IN_from_sum[13][60] , \ADDER_IN_from_sum[13][59] , 
        \ADDER_IN_from_sum[13][58] , \ADDER_IN_from_sum[13][57] , 
        \ADDER_IN_from_sum[13][56] , \ADDER_IN_from_sum[13][55] , 
        \ADDER_IN_from_sum[13][54] , \ADDER_IN_from_sum[13][53] , 
        \ADDER_IN_from_sum[13][52] , \ADDER_IN_from_sum[13][51] , 
        \ADDER_IN_from_sum[13][50] , \ADDER_IN_from_sum[13][49] , 
        \ADDER_IN_from_sum[13][48] , \ADDER_IN_from_sum[13][47] , 
        \ADDER_IN_from_sum[13][46] , \ADDER_IN_from_sum[13][45] , 
        \ADDER_IN_from_sum[13][44] , \ADDER_IN_from_sum[13][43] , 
        \ADDER_IN_from_sum[13][42] , \ADDER_IN_from_sum[13][41] , 
        \ADDER_IN_from_sum[13][40] , \ADDER_IN_from_sum[13][39] , 
        \ADDER_IN_from_sum[13][38] , \ADDER_IN_from_sum[13][37] , 
        \ADDER_IN_from_sum[13][36] , \ADDER_IN_from_sum[13][35] , 
        \ADDER_IN_from_sum[13][34] , \ADDER_IN_from_sum[13][33] , 
        \ADDER_IN_from_sum[13][32] , \ADDER_IN_from_sum[13][31] , 
        \ADDER_IN_from_sum[13][30] , \ADDER_IN_from_sum[13][29] , 
        \ADDER_IN_from_sum[13][28] , \ADDER_IN_from_sum[13][27] , 
        \ADDER_IN_from_sum[13][26] , \ADDER_IN_from_sum[13][25] , 
        \ADDER_IN_from_sum[13][24] , \ADDER_IN_from_sum[13][23] , 
        \ADDER_IN_from_sum[13][22] , \ADDER_IN_from_sum[13][21] , 
        \ADDER_IN_from_sum[13][20] , \ADDER_IN_from_sum[13][19] , 
        \ADDER_IN_from_sum[13][18] , \ADDER_IN_from_sum[13][17] , 
        \ADDER_IN_from_sum[13][16] , \ADDER_IN_from_sum[13][15] , 
        \ADDER_IN_from_sum[13][14] , \ADDER_IN_from_sum[13][13] , 
        \ADDER_IN_from_sum[13][12] , \ADDER_IN_from_sum[13][11] , 
        \ADDER_IN_from_sum[13][10] , \ADDER_IN_from_sum[13][9] , 
        \ADDER_IN_from_sum[13][8] , \ADDER_IN_from_sum[13][7] , 
        \ADDER_IN_from_sum[13][6] , \ADDER_IN_from_sum[13][5] , 
        \ADDER_IN_from_sum[13][4] , \ADDER_IN_from_sum[13][3] , 
        \ADDER_IN_from_sum[13][2] , \ADDER_IN_from_sum[13][1] , 
        \ADDER_IN_from_sum[13][0] }), .B({\ADDER_IN_from_mux[15][63] , 
        \ADDER_IN_from_mux[15][62] , \ADDER_IN_from_mux[15][61] , 
        \ADDER_IN_from_mux[15][60] , \ADDER_IN_from_mux[15][59] , 
        \ADDER_IN_from_mux[15][58] , \ADDER_IN_from_mux[15][57] , 
        \ADDER_IN_from_mux[15][56] , \ADDER_IN_from_mux[15][55] , 
        \ADDER_IN_from_mux[15][54] , \ADDER_IN_from_mux[15][53] , 
        \ADDER_IN_from_mux[15][52] , \ADDER_IN_from_mux[15][51] , 
        \ADDER_IN_from_mux[15][50] , \ADDER_IN_from_mux[15][49] , 
        \ADDER_IN_from_mux[15][48] , \ADDER_IN_from_mux[15][47] , 
        \ADDER_IN_from_mux[15][46] , \ADDER_IN_from_mux[15][45] , 
        \ADDER_IN_from_mux[15][44] , \ADDER_IN_from_mux[15][43] , 
        \ADDER_IN_from_mux[15][42] , \ADDER_IN_from_mux[15][41] , 
        \ADDER_IN_from_mux[15][40] , \ADDER_IN_from_mux[15][39] , 
        \ADDER_IN_from_mux[15][38] , \ADDER_IN_from_mux[15][37] , 
        \ADDER_IN_from_mux[15][36] , \ADDER_IN_from_mux[15][35] , 
        \ADDER_IN_from_mux[15][34] , \ADDER_IN_from_mux[15][33] , 
        \ADDER_IN_from_mux[15][32] , \ADDER_IN_from_mux[15][31] , 
        \ADDER_IN_from_mux[15][30] , \ADDER_IN_from_mux[15][29] , 
        \ADDER_IN_from_mux[15][28] , \ADDER_IN_from_mux[15][27] , 
        \ADDER_IN_from_mux[15][26] , \ADDER_IN_from_mux[15][25] , 
        \ADDER_IN_from_mux[15][24] , \ADDER_IN_from_mux[15][23] , 
        \ADDER_IN_from_mux[15][22] , \ADDER_IN_from_mux[15][21] , 
        \ADDER_IN_from_mux[15][20] , \ADDER_IN_from_mux[15][19] , 
        \ADDER_IN_from_mux[15][18] , \ADDER_IN_from_mux[15][17] , 
        \ADDER_IN_from_mux[15][16] , \ADDER_IN_from_mux[15][15] , 
        \ADDER_IN_from_mux[15][14] , \ADDER_IN_from_mux[15][13] , 
        \ADDER_IN_from_mux[15][12] , \ADDER_IN_from_mux[15][11] , 
        \ADDER_IN_from_mux[15][10] , \ADDER_IN_from_mux[15][9] , 
        \ADDER_IN_from_mux[15][8] , \ADDER_IN_from_mux[15][7] , 
        \ADDER_IN_from_mux[15][6] , \ADDER_IN_from_mux[15][5] , 
        \ADDER_IN_from_mux[15][4] , \ADDER_IN_from_mux[15][3] , 
        \ADDER_IN_from_mux[15][2] , \ADDER_IN_from_mux[15][1] , 
        \ADDER_IN_from_mux[15][0] }), .S({\ADDER_IN_from_sum[14][63] , 
        \ADDER_IN_from_sum[14][62] , \ADDER_IN_from_sum[14][61] , 
        \ADDER_IN_from_sum[14][60] , \ADDER_IN_from_sum[14][59] , 
        \ADDER_IN_from_sum[14][58] , \ADDER_IN_from_sum[14][57] , 
        \ADDER_IN_from_sum[14][56] , \ADDER_IN_from_sum[14][55] , 
        \ADDER_IN_from_sum[14][54] , \ADDER_IN_from_sum[14][53] , 
        \ADDER_IN_from_sum[14][52] , \ADDER_IN_from_sum[14][51] , 
        \ADDER_IN_from_sum[14][50] , \ADDER_IN_from_sum[14][49] , 
        \ADDER_IN_from_sum[14][48] , \ADDER_IN_from_sum[14][47] , 
        \ADDER_IN_from_sum[14][46] , \ADDER_IN_from_sum[14][45] , 
        \ADDER_IN_from_sum[14][44] , \ADDER_IN_from_sum[14][43] , 
        \ADDER_IN_from_sum[14][42] , \ADDER_IN_from_sum[14][41] , 
        \ADDER_IN_from_sum[14][40] , \ADDER_IN_from_sum[14][39] , 
        \ADDER_IN_from_sum[14][38] , \ADDER_IN_from_sum[14][37] , 
        \ADDER_IN_from_sum[14][36] , \ADDER_IN_from_sum[14][35] , 
        \ADDER_IN_from_sum[14][34] , \ADDER_IN_from_sum[14][33] , 
        \ADDER_IN_from_sum[14][32] , \ADDER_IN_from_sum[14][31] , 
        \ADDER_IN_from_sum[14][30] , \ADDER_IN_from_sum[14][29] , 
        \ADDER_IN_from_sum[14][28] , \ADDER_IN_from_sum[14][27] , 
        \ADDER_IN_from_sum[14][26] , \ADDER_IN_from_sum[14][25] , 
        \ADDER_IN_from_sum[14][24] , \ADDER_IN_from_sum[14][23] , 
        \ADDER_IN_from_sum[14][22] , \ADDER_IN_from_sum[14][21] , 
        \ADDER_IN_from_sum[14][20] , \ADDER_IN_from_sum[14][19] , 
        \ADDER_IN_from_sum[14][18] , \ADDER_IN_from_sum[14][17] , 
        \ADDER_IN_from_sum[14][16] , \ADDER_IN_from_sum[14][15] , 
        \ADDER_IN_from_sum[14][14] , \ADDER_IN_from_sum[14][13] , 
        \ADDER_IN_from_sum[14][12] , \ADDER_IN_from_sum[14][11] , 
        \ADDER_IN_from_sum[14][10] , \ADDER_IN_from_sum[14][9] , 
        \ADDER_IN_from_sum[14][8] , \ADDER_IN_from_sum[14][7] , 
        \ADDER_IN_from_sum[14][6] , \ADDER_IN_from_sum[14][5] , 
        \ADDER_IN_from_sum[14][4] , \ADDER_IN_from_sum[14][3] , 
        \ADDER_IN_from_sum[14][2] , \ADDER_IN_from_sum[14][1] , 
        \ADDER_IN_from_sum[14][0] }) );
  FD_GENERIC_NBIT64 reg_out ( .D({\ADDER_IN_from_sum[14][63] , 
        \ADDER_IN_from_sum[14][62] , \ADDER_IN_from_sum[14][61] , 
        \ADDER_IN_from_sum[14][60] , \ADDER_IN_from_sum[14][59] , 
        \ADDER_IN_from_sum[14][58] , \ADDER_IN_from_sum[14][57] , 
        \ADDER_IN_from_sum[14][56] , \ADDER_IN_from_sum[14][55] , 
        \ADDER_IN_from_sum[14][54] , \ADDER_IN_from_sum[14][53] , 
        \ADDER_IN_from_sum[14][52] , \ADDER_IN_from_sum[14][51] , 
        \ADDER_IN_from_sum[14][50] , \ADDER_IN_from_sum[14][49] , 
        \ADDER_IN_from_sum[14][48] , \ADDER_IN_from_sum[14][47] , 
        \ADDER_IN_from_sum[14][46] , \ADDER_IN_from_sum[14][45] , 
        \ADDER_IN_from_sum[14][44] , \ADDER_IN_from_sum[14][43] , 
        \ADDER_IN_from_sum[14][42] , \ADDER_IN_from_sum[14][41] , 
        \ADDER_IN_from_sum[14][40] , \ADDER_IN_from_sum[14][39] , 
        \ADDER_IN_from_sum[14][38] , \ADDER_IN_from_sum[14][37] , 
        \ADDER_IN_from_sum[14][36] , \ADDER_IN_from_sum[14][35] , 
        \ADDER_IN_from_sum[14][34] , \ADDER_IN_from_sum[14][33] , 
        \ADDER_IN_from_sum[14][32] , \ADDER_IN_from_sum[14][31] , 
        \ADDER_IN_from_sum[14][30] , \ADDER_IN_from_sum[14][29] , 
        \ADDER_IN_from_sum[14][28] , \ADDER_IN_from_sum[14][27] , 
        \ADDER_IN_from_sum[14][26] , \ADDER_IN_from_sum[14][25] , 
        \ADDER_IN_from_sum[14][24] , \ADDER_IN_from_sum[14][23] , 
        \ADDER_IN_from_sum[14][22] , \ADDER_IN_from_sum[14][21] , 
        \ADDER_IN_from_sum[14][20] , \ADDER_IN_from_sum[14][19] , 
        \ADDER_IN_from_sum[14][18] , \ADDER_IN_from_sum[14][17] , 
        \ADDER_IN_from_sum[14][16] , \ADDER_IN_from_sum[14][15] , 
        \ADDER_IN_from_sum[14][14] , \ADDER_IN_from_sum[14][13] , 
        \ADDER_IN_from_sum[14][12] , \ADDER_IN_from_sum[14][11] , 
        \ADDER_IN_from_sum[14][10] , \ADDER_IN_from_sum[14][9] , 
        \ADDER_IN_from_sum[14][8] , \ADDER_IN_from_sum[14][7] , 
        \ADDER_IN_from_sum[14][6] , \ADDER_IN_from_sum[14][5] , 
        \ADDER_IN_from_sum[14][4] , \ADDER_IN_from_sum[14][3] , 
        \ADDER_IN_from_sum[14][2] , \ADDER_IN_from_sum[14][1] , 
        \ADDER_IN_from_sum[14][0] }), .CLK(Clk), .RESET(reset), .Q(MUL_OUT) );
  BUF_X1 U2 ( .A(in_1[9]), .Z(n539) );
  BUF_X1 U3 ( .A(in_1[8]), .Z(n536) );
  BUF_X1 U4 ( .A(in_1[7]), .Z(n533) );
  BUF_X1 U5 ( .A(in_1[0]), .Z(n511) );
  BUF_X1 U6 ( .A(in_1[17]), .Z(n568) );
  BUF_X2 U7 ( .A(in_1[14]), .Z(n555) );
  BUF_X1 U8 ( .A(n577), .Z(n580) );
  BUF_X1 U9 ( .A(n577), .Z(n579) );
  BUF_X2 U10 ( .A(in_1[12]), .Z(n551) );
  BUF_X4 U11 ( .A(in_1[7]), .Z(n531) );
  BUF_X1 U12 ( .A(n511), .Z(n510) );
  CLKBUF_X2 U13 ( .A(in_1[6]), .Z(n530) );
  CLKBUF_X2 U14 ( .A(n519), .Z(n521) );
  BUF_X2 U15 ( .A(n511), .Z(n509) );
  INV_X2 U16 ( .A(n492), .ZN(n493) );
  BUF_X2 U17 ( .A(n517), .Z(n504) );
  BUF_X2 U18 ( .A(n525), .Z(n490) );
  CLKBUF_X1 U19 ( .A(in_1[5]), .Z(n525) );
  BUF_X4 U20 ( .A(n529), .Z(n491) );
  INV_X1 U21 ( .A(n509), .ZN(n492) );
  BUF_X2 U22 ( .A(in_1[3]), .Z(n494) );
  CLKBUF_X1 U23 ( .A(in_1[3]), .Z(n495) );
  BUF_X1 U24 ( .A(in_1[3]), .Z(n520) );
  BUF_X1 U25 ( .A(n526), .Z(n501) );
  BUF_X2 U26 ( .A(n524), .Z(n528) );
  CLKBUF_X1 U27 ( .A(n543), .Z(n546) );
  CLKBUF_X2 U28 ( .A(n510), .Z(n507) );
  CLKBUF_X1 U29 ( .A(in_1[0]), .Z(n497) );
  BUF_X1 U30 ( .A(n524), .Z(n526) );
  BUF_X1 U31 ( .A(in_1[5]), .Z(n524) );
  BUF_X1 U32 ( .A(in_1[4]), .Z(n505) );
  CLKBUF_X1 U33 ( .A(in_1[4]), .Z(n523) );
  CLKBUF_X1 U34 ( .A(in_1[4]), .Z(n522) );
  CLKBUF_X1 U35 ( .A(in_1[3]), .Z(n519) );
  BUF_X4 U36 ( .A(in_1[9]), .Z(n538) );
  CLKBUF_X1 U37 ( .A(in_1[9]), .Z(n537) );
  BUF_X2 U38 ( .A(n523), .Z(n496) );
  BUF_X2 U39 ( .A(n516), .Z(n517) );
  BUF_X2 U40 ( .A(in_1[2]), .Z(n516) );
  CLKBUF_X1 U41 ( .A(n516), .Z(n518) );
  BUF_X2 U42 ( .A(n558), .Z(n562) );
  BUF_X2 U43 ( .A(n584), .Z(n586) );
  CLKBUF_X2 U44 ( .A(in_1[16]), .Z(n565) );
  CLKBUF_X1 U45 ( .A(n511), .Z(n498) );
  BUF_X2 U46 ( .A(n685), .Z(n654) );
  BUF_X2 U47 ( .A(n690), .Z(n641) );
  BUF_X2 U48 ( .A(n685), .Z(n655) );
  BUF_X2 U49 ( .A(n689), .Z(n642) );
  BUF_X2 U50 ( .A(n686), .Z(n652) );
  BUF_X2 U51 ( .A(n688), .Z(n647) );
  BUF_X2 U52 ( .A(n689), .Z(n644) );
  BUF_X2 U53 ( .A(n687), .Z(n649) );
  BUF_X2 U54 ( .A(n687), .Z(n648) );
  BUF_X2 U55 ( .A(n689), .Z(n643) );
  BUF_X2 U56 ( .A(n691), .Z(n638) );
  BUF_X2 U57 ( .A(n690), .Z(n640) );
  BUF_X2 U58 ( .A(n690), .Z(n639) );
  BUF_X2 U59 ( .A(n691), .Z(n637) );
  BUF_X2 U60 ( .A(n691), .Z(n636) );
  CLKBUF_X1 U61 ( .A(n558), .Z(n560) );
  BUF_X2 U62 ( .A(n578), .Z(n583) );
  CLKBUF_X1 U63 ( .A(n558), .Z(n561) );
  BUF_X4 U64 ( .A(n543), .Z(n545) );
  BUF_X4 U65 ( .A(n569), .Z(n572) );
  BUF_X4 U66 ( .A(n512), .Z(n515) );
  BUF_X4 U67 ( .A(n590), .Z(n593) );
  CLKBUF_X1 U68 ( .A(n569), .Z(n573) );
  BUF_X2 U69 ( .A(in_1[28]), .Z(n617) );
  BUF_X2 U70 ( .A(in_1[30]), .Z(n626) );
  BUF_X2 U71 ( .A(in_1[26]), .Z(n611) );
  BUF_X2 U72 ( .A(in_1[22]), .Z(n596) );
  BUF_X2 U73 ( .A(in_1[18]), .Z(n574) );
  BUF_X2 U74 ( .A(in_1[25]), .Z(n608) );
  BUF_X2 U75 ( .A(in_1[12]), .Z(n549) );
  BUF_X2 U76 ( .A(in_1[8]), .Z(n534) );
  CLKBUF_X1 U77 ( .A(in_1[15]), .Z(n559) );
  BUF_X2 U78 ( .A(in_1[1]), .Z(n512) );
  CLKBUF_X3 U79 ( .A(n686), .Z(n653) );
  BUF_X2 U80 ( .A(n686), .Z(n651) );
  BUF_X2 U81 ( .A(n682), .Z(n664) );
  BUF_X2 U82 ( .A(n679), .Z(n672) );
  BUF_X2 U83 ( .A(n680), .Z(n671) );
  BUF_X2 U84 ( .A(n682), .Z(n663) );
  BUF_X2 U85 ( .A(n679), .Z(n673) );
  BUF_X2 U86 ( .A(n684), .Z(n658) );
  CLKBUF_X3 U87 ( .A(n679), .Z(n674) );
  BUF_X2 U88 ( .A(n684), .Z(n657) );
  BUF_X2 U89 ( .A(n684), .Z(n659) );
  BUF_X1 U90 ( .A(n678), .Z(n677) );
  BUF_X2 U91 ( .A(n688), .Z(n646) );
  BUF_X2 U92 ( .A(n688), .Z(n645) );
  BUF_X2 U93 ( .A(n687), .Z(n650) );
  BUF_X2 U94 ( .A(n685), .Z(n656) );
  BUF_X2 U95 ( .A(n682), .Z(n665) );
  BUF_X2 U96 ( .A(n680), .Z(n669) );
  BUF_X2 U97 ( .A(n681), .Z(n667) );
  BUF_X2 U98 ( .A(n681), .Z(n668) );
  CLKBUF_X3 U99 ( .A(n678), .Z(n675) );
  CLKBUF_X3 U100 ( .A(n678), .Z(n676) );
  BUF_X2 U101 ( .A(n683), .Z(n660) );
  BUF_X2 U102 ( .A(n683), .Z(n661) );
  BUF_X2 U103 ( .A(n680), .Z(n670) );
  BUF_X2 U104 ( .A(n681), .Z(n666) );
  BUF_X2 U105 ( .A(n683), .Z(n662) );
  CLKBUF_X1 U106 ( .A(n494), .Z(n499) );
  CLKBUF_X1 U107 ( .A(n517), .Z(n503) );
  CLKBUF_X1 U108 ( .A(n494), .Z(n500) );
  BUF_X1 U109 ( .A(n632), .Z(n687) );
  BUF_X1 U110 ( .A(n632), .Z(n689) );
  BUF_X1 U111 ( .A(n631), .Z(n685) );
  BUF_X1 U112 ( .A(n632), .Z(n688) );
  BUF_X1 U113 ( .A(n631), .Z(n686) );
  BUF_X1 U114 ( .A(n629), .Z(n680) );
  BUF_X1 U115 ( .A(n629), .Z(n679) );
  BUF_X1 U116 ( .A(n630), .Z(n682) );
  BUF_X1 U117 ( .A(n631), .Z(n684) );
  BUF_X1 U118 ( .A(n633), .Z(n690) );
  BUF_X1 U119 ( .A(n629), .Z(n678) );
  BUF_X1 U120 ( .A(n630), .Z(n681) );
  BUF_X1 U121 ( .A(n633), .Z(n691) );
  BUF_X1 U122 ( .A(n630), .Z(n683) );
  BUF_X2 U123 ( .A(n512), .Z(n513) );
  BUF_X1 U124 ( .A(n577), .Z(n581) );
  BUF_X2 U125 ( .A(n512), .Z(n514) );
  BUF_X1 U126 ( .A(n559), .Z(n563) );
  BUF_X1 U127 ( .A(n559), .Z(n564) );
  BUF_X4 U128 ( .A(n568), .Z(n570) );
  BUF_X1 U129 ( .A(n578), .Z(n582) );
  BUF_X2 U130 ( .A(n602), .Z(n605) );
  BUF_X2 U131 ( .A(n590), .Z(n592) );
  BUF_X2 U132 ( .A(n602), .Z(n604) );
  BUF_X4 U133 ( .A(n568), .Z(n571) );
  BUF_X2 U134 ( .A(n584), .Z(n587) );
  BUF_X2 U135 ( .A(n620), .Z(n622) );
  BUF_X2 U136 ( .A(n591), .Z(n594) );
  BUF_X2 U137 ( .A(n620), .Z(n623) );
  BUF_X2 U138 ( .A(n603), .Z(n606) );
  BUF_X2 U139 ( .A(n585), .Z(n588) );
  BUF_X2 U140 ( .A(n621), .Z(n624) );
  BUF_X2 U141 ( .A(n544), .Z(n547) );
  BUF_X2 U142 ( .A(n524), .Z(n527) );
  BUF_X1 U143 ( .A(n621), .Z(n625) );
  BUF_X1 U144 ( .A(n544), .Z(n548) );
  BUF_X1 U145 ( .A(n603), .Z(n607) );
  BUF_X1 U146 ( .A(n591), .Z(n595) );
  BUF_X1 U147 ( .A(n585), .Z(n589) );
  BUF_X1 U148 ( .A(n634), .Z(n632) );
  BUF_X1 U149 ( .A(n634), .Z(n631) );
  BUF_X1 U150 ( .A(n635), .Z(n630) );
  BUF_X1 U151 ( .A(n635), .Z(n629) );
  BUF_X1 U152 ( .A(n634), .Z(n633) );
  BUF_X2 U153 ( .A(in_1[28]), .Z(n619) );
  BUF_X2 U154 ( .A(in_1[22]), .Z(n598) );
  BUF_X4 U155 ( .A(in_1[13]), .Z(n552) );
  BUF_X4 U156 ( .A(in_1[10]), .Z(n540) );
  BUF_X4 U157 ( .A(in_1[18]), .Z(n575) );
  BUF_X4 U158 ( .A(in_1[10]), .Z(n541) );
  BUF_X1 U159 ( .A(in_1[30]), .Z(n628) );
  BUF_X2 U160 ( .A(in_1[28]), .Z(n618) );
  BUF_X4 U161 ( .A(in_1[6]), .Z(n529) );
  BUF_X4 U162 ( .A(in_1[22]), .Z(n597) );
  BUF_X4 U163 ( .A(in_1[14]), .Z(n556) );
  BUF_X4 U164 ( .A(in_1[12]), .Z(n550) );
  BUF_X2 U165 ( .A(in_1[30]), .Z(n627) );
  BUF_X4 U166 ( .A(in_1[13]), .Z(n553) );
  BUF_X4 U167 ( .A(in_1[26]), .Z(n612) );
  BUF_X2 U168 ( .A(in_1[23]), .Z(n599) );
  BUF_X2 U169 ( .A(in_1[27]), .Z(n614) );
  BUF_X4 U170 ( .A(in_1[8]), .Z(n535) );
  BUF_X4 U171 ( .A(in_1[7]), .Z(n532) );
  BUF_X4 U172 ( .A(in_1[23]), .Z(n600) );
  BUF_X4 U173 ( .A(in_1[16]), .Z(n566) );
  BUF_X2 U174 ( .A(in_1[27]), .Z(n615) );
  BUF_X4 U175 ( .A(in_1[25]), .Z(n609) );
  BUF_X1 U176 ( .A(in_1[24]), .Z(n602) );
  BUF_X1 U177 ( .A(in_1[21]), .Z(n590) );
  BUF_X1 U178 ( .A(in_1[20]), .Z(n584) );
  BUF_X1 U179 ( .A(in_1[11]), .Z(n543) );
  BUF_X1 U180 ( .A(in_1[29]), .Z(n620) );
  CLKBUF_X1 U181 ( .A(in_1[11]), .Z(n544) );
  BUF_X1 U182 ( .A(in_1[29]), .Z(n621) );
  BUF_X1 U183 ( .A(in_1[17]), .Z(n569) );
  CLKBUF_X1 U184 ( .A(in_1[20]), .Z(n585) );
  CLKBUF_X1 U185 ( .A(in_1[21]), .Z(n591) );
  BUF_X1 U186 ( .A(in_1[24]), .Z(n603) );
  BUF_X1 U187 ( .A(in_1[19]), .Z(n578) );
  CLKBUF_X1 U188 ( .A(in_1[19]), .Z(n577) );
  BUF_X1 U189 ( .A(in_1[15]), .Z(n558) );
  BUF_X1 U190 ( .A(in_1[31]), .Z(n634) );
  BUF_X1 U191 ( .A(in_1[31]), .Z(n635) );
  BUF_X1 U192 ( .A(n516), .Z(n502) );
  BUF_X4 U193 ( .A(in_1[4]), .Z(n506) );
  CLKBUF_X1 U194 ( .A(n511), .Z(n508) );
  BUF_X4 U195 ( .A(in_1[10]), .Z(n542) );
  BUF_X4 U196 ( .A(in_1[13]), .Z(n554) );
  BUF_X4 U197 ( .A(in_1[14]), .Z(n557) );
  BUF_X4 U198 ( .A(in_1[16]), .Z(n567) );
  BUF_X4 U199 ( .A(in_1[18]), .Z(n576) );
  BUF_X4 U200 ( .A(in_1[23]), .Z(n601) );
  BUF_X4 U201 ( .A(in_1[25]), .Z(n610) );
  BUF_X4 U202 ( .A(in_1[26]), .Z(n613) );
  BUF_X4 U203 ( .A(in_1[27]), .Z(n616) );
endmodule

